CNP Edge Only Rom		"0", "1", "2", "3", "4", "5", "20", "21", "22", "23", "24", "25", "26", "27", "28", "29", "30", "31", "39", "40", "41", "42", "43", "44", "45", "46", "47", "48", "49", "50", "58", "59", "60", "61", "62", "63", "64", "65", "66", "67", "68", "69", "70", "71", "72", "73", "74", "75", "6", "7", "8", "9", "10", "11", "12", "13", "14", "15", "16", "17", "18", "19", "32", "33", "34", "35", "36", "37", "38", "51", "52", "53", "54", "55", "56", "57", 
CNP Edge+Restart Rom	"0", "1", "2", "3", "4", "133", "20", "21", "22", "23", "24", "153", "26", "27", "28", "29", "30", "159", "39", "40", "41", "42", "43", "172", "45", "46", "47", "48", "49", "178", "58", "59", "60", "61", "62", "191", "64", "65", "66", "67", "68", "197", "70", "71", "72", "73", "74", "203", "6", "7", "8", "9", "10", "11", "140", "13", "14", "15", "16", "17", "18", "147", "32", "33", "34", "35", "36", "37", "166", "51", "52", "53", "54", "55", "56", "185", 
CNP Rotation Rom		"2", "23", "41", "13", "89", "96", "35", "49", "31", "71", "96", "96", "57", "12", "55", "24", "96", "96", "1", "43", "82", "78", "96", "96", "85", "23", "94", "49", "96", "96", "2", "37", "26", "24", "96", "96", "89", "31", "57", "47", "96", "96", "53", "30", "55", "70", "89", "96", "69", "74", "17", "87", "84", "96", "96", "72", "74", "15", "63", "96", "96", "96", "50", "56", "14", "17", "96", "96", "96", "84", "13", "72", "53", "45", "96", "96", 


VNP Edge Only Rom		5, 11, 89, 12, 18, 90, 19, 24, 91, 25, 30, 92, 31, 37, 93, 38, 43, 94, 44, 49, 95, 50, 56, 96, 57, 62, 97, 63, 68, 98, 69, 75, 99, 20, 51, 70, 76, 0, 6, 45, 77, 13, 40, 65, 79, 14, 32, 52, 80, 8, 27, 47, 82, 2, 22, 66, 84, 29, 42, 60, 86, 4, 36, 74, 88, 1, 21, 26, 39, 46, 64, 78, 7, 15, 33, 53, 58, 71, 81, 9, 16, 34, 54, 59, 72, 83, 3, 23, 28, 41, 48, 67, 85, 10, 17, 35, 55, 61, 73, 87, 
VNP Edge+Restart Rom	"00000101", "00001011", "11011001", "00001100", "00010010", "11011010", "00010011", "00011000", "11011011", "00011001", "00011110", "11011100", "00011111", "00100101", "11011101", "00100110", "00101011", "11011110", "00101100", "00110001", "11011111", "00110010", "00111000", "11100000", "00111001", "00111110", "11100001", "00111111", "01000100", "11100010", "01000101", "01001011", "11100011", "00010100", "00110011", "01000110", "11001100", "00000000", "00000110", "00101101", "11001101", "00001101", "00101000", "01000001", "11001111", "00001110", "00100000", "00110100", "11010000", "00001000", "00011011", "00101111", "11010010", "00000010", "00010110", "01000010", "11010100", "00011101", "00101010", "00111100", "11010110", "00000100", "00100100", "01001010", "11011000", "00000001", "00010101", "00011010", "00100111", "00101110", "01000000", "11001110", "00000111", "00001111", "00100001", "00110101", "00111010", "01000111", "11010001", "00001001", "00010000", "00100010", "00110110", "00111011", "01001000", "11010011", "00000011", "00010111", "00011100", "00101001", "00110000", "01000011", "11010101", "00001010", "00010001", "00100011", "00110111", "00111101", "01001001", "11010111", 
VNP Rotation Rom		0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 12, 43, 0, 94, 27, 11, 0, 24, 53, 65, 0, 22, 46, 83, 0, 79, 84, 2, 0, 55, 65, 39, 0, 72, 18, 70, 0, 7, 0, 7, 0, 73, 47, 39, 95, 73, 7, 0, 22, 81, 40, 24, 94, 66, 0, 9, 33, 82, 43, 59, 41, 0, 83, 25, 41, 14, 47, 49, 0, 12, 0, 79, 51, 72, 26, 0, 
