LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CNP_Input_Edge_Memory is
	Port (
		clk			: in  std_logic;

		RdAddr		: in  std_logic_vector(13 downto 0);
		Do			: out std_logic_vector(11 downto 0)
	);
end CNP_Input_Edge_Memory;

architecture Behavioral of CNP_Input_Edge_Memory is
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 11672-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
24,   25,   26+2048
,   51,   52,   53+2048
,   54,   55,   56+2048
,   57,   58,   59+2048
,   76,   77,   78+2048
,   99,  100,  101+2048
,  102,  103,  104+2048
,  105,  106,  107+2048
,  112,  113,  114+2048
,  159,  160,  161+2048
,  186,  187,  188+2048
,  189,  190,  191+2048
,  192,  193,  194+2048
,  211,  212,  213+2048
,  234,  235,  236+2048
,  237,  238,  239+2048
,  240,  241,  242+2048
,  247,  248,  249+2048
,  294,  295,  296+2048
,  321,  322,  323+2048
,  324,  325,  326+2048
,  327,  328,  329+2048
,  346,  347,  348+2048
,  369,  370,  371+2048
,  372,  373,  374+2048
,  375,  376,  377+2048
,  382,  383,  384+2048
,  429,  430,  431+2048
,  456,  457,  458+2048
,  459,  460,  461+2048
,  462,  463,  464+2048
,  481,  482,  483+2048
,  504,  505,  506+2048
,  507,  508,  509+2048
,  510,  511,  512+2048
,  517,  518,  519+2048
,  564,  565,  566+2048
,  591,  592,  593+2048
,  594,  595,  596+2048
,  597,  598,  599+2048
,  616,  617,  618+2048
,  639,  640,  641+2048
,  642,  643,  644+2048
,  645,  646,  647+2048
,  652,  653,  654+2048
,  699,  700,  701+2048
,  726,  727,  728+2048
,  729,  730,  731+2048
,  732,  733,  734+2048
,  751,  752,  753+2048
,  774,  775,  776+2048
,  777,  778,  779+2048
,  780,  781,  782+2048
,  787,  788,  789+2048
,  834,  835,  836+2048
,  861,  862,  863+2048
,  864,  865,  866+2048
,  867,  868,  869+2048
,  886,  887,  888+2048
,  909,  910,  911+2048
,  912,  913,  914+2048
,  915,  916,  917+2048
,  922,  923,  924+2048
,  969,  970,  971+2048
,  996,  997,  998+2048
,  999, 1000, 1001+2048
, 1002, 1003, 1004+2048
, 1021, 1022, 1023+2048
, 1044, 1045, 1046+2048
, 1047, 1048, 1049+2048
, 1050, 1051, 1052+2048
, 1057, 1058, 1059+2048
,    0,    1,    2,    3+2048
,    4,    5,    6,    7+2048
,    8,    9,   10,   11+2048
,   12,   13,   14,   15+2048
,   16,   17,   18,   19+2048
,   20,   21,   22,   23+2048
,   27,   28,   29,   30+2048
,   31,   32,   33,   34+2048
,   35,   36,   37,   38+2048
,   39,   40,   41,   42+2048
,   43,   44,   45,   46+2048
,   47,   48,   49,   50+2048
,   60,   61,   62,   63+2048
,   64,   65,   66,   67+2048
,   68,   69,   70,   71+2048
,   72,   73,   74,   75+2048
,   79,   80,   81,   82+2048
,   83,   84,   85,   86+2048
,   87,   88,   89,   90+2048
,   91,   92,   93,   94+2048
,   95,   96,   97,   98+2048
,  108,  109,  110,  111+2048
,  115,  116,  117,  118+2048
,  119,  120,  121,  122+2048
,  123,  124,  125,  126+2048
,  127,  128,  129,  130+2048
,  131,  132,  133,  134+2048
,  135,  136,  137,  138+2048
,  139,  140,  141,  142+2048
,  143,  144,  145,  146+2048
,  147,  148,  149,  150+2048
,  151,  152,  153,  154+2048
,  155,  156,  157,  158+2048
,  162,  163,  164,  165+2048
,  166,  167,  168,  169+2048
,  170,  171,  172,  173+2048
,  174,  175,  176,  177+2048
,  178,  179,  180,  181+2048
,  182,  183,  184,  185+2048
,  195,  196,  197,  198+2048
,  199,  200,  201,  202+2048
,  203,  204,  205,  206+2048
,  207,  208,  209,  210+2048
,  214,  215,  216,  217+2048
,  218,  219,  220,  221+2048
,  222,  223,  224,  225+2048
,  226,  227,  228,  229+2048
,  230,  231,  232,  233+2048
,  243,  244,  245,  246+2048
,  250,  251,  252,  253+2048
,  254,  255,  256,  257+2048
,  258,  259,  260,  261+2048
,  262,  263,  264,  265+2048
,  266,  267,  268,  269+2048
,  270,  271,  272,  273+2048
,  274,  275,  276,  277+2048
,  278,  279,  280,  281+2048
,  282,  283,  284,  285+2048
,  286,  287,  288,  289+2048
,  290,  291,  292,  293+2048
,  297,  298,  299,  300+2048
,  301,  302,  303,  304+2048
,  305,  306,  307,  308+2048
,  309,  310,  311,  312+2048
,  313,  314,  315,  316+2048
,  317,  318,  319,  320+2048
,  330,  331,  332,  333+2048
,  334,  335,  336,  337+2048
,  338,  339,  340,  341+2048
,  342,  343,  344,  345+2048
,  349,  350,  351,  352+2048
,  353,  354,  355,  356+2048
,  357,  358,  359,  360+2048
,  361,  362,  363,  364+2048
,  365,  366,  367,  368+2048
,  378,  379,  380,  381+2048
,  385,  386,  387,  388+2048
,  389,  390,  391,  392+2048
,  393,  394,  395,  396+2048
,  397,  398,  399,  400+2048
,  401,  402,  403,  404+2048
,  405,  406,  407,  408+2048
,  409,  410,  411,  412+2048
,  413,  414,  415,  416+2048
,  417,  418,  419,  420+2048
,  421,  422,  423,  424+2048
,  425,  426,  427,  428+2048
,  432,  433,  434,  435+2048
,  436,  437,  438,  439+2048
,  440,  441,  442,  443+2048
,  444,  445,  446,  447+2048
,  448,  449,  450,  451+2048
,  452,  453,  454,  455+2048
,  465,  466,  467,  468+2048
,  469,  470,  471,  472+2048
,  473,  474,  475,  476+2048
,  477,  478,  479,  480+2048
,  484,  485,  486,  487+2048
,  488,  489,  490,  491+2048
,  492,  493,  494,  495+2048
,  496,  497,  498,  499+2048
,  500,  501,  502,  503+2048
,  513,  514,  515,  516+2048
,  520,  521,  522,  523+2048
,  524,  525,  526,  527+2048
,  528,  529,  530,  531+2048
,  532,  533,  534,  535+2048
,  536,  537,  538,  539+2048
,  540,  541,  542,  543+2048
,  544,  545,  546,  547+2048
,  548,  549,  550,  551+2048
,  552,  553,  554,  555+2048
,  556,  557,  558,  559+2048
,  560,  561,  562,  563+2048
,  567,  568,  569,  570+2048
,  571,  572,  573,  574+2048
,  575,  576,  577,  578+2048
,  579,  580,  581,  582+2048
,  583,  584,  585,  586+2048
,  587,  588,  589,  590+2048
,  600,  601,  602,  603+2048
,  604,  605,  606,  607+2048
,  608,  609,  610,  611+2048
,  612,  613,  614,  615+2048
,  619,  620,  621,  622+2048
,  623,  624,  625,  626+2048
,  627,  628,  629,  630+2048
,  631,  632,  633,  634+2048
,  635,  636,  637,  638+2048
,  648,  649,  650,  651+2048
,  655,  656,  657,  658+2048
,  659,  660,  661,  662+2048
,  663,  664,  665,  666+2048
,  667,  668,  669,  670+2048
,  671,  672,  673,  674+2048
,  675,  676,  677,  678+2048
,  679,  680,  681,  682+2048
,  683,  684,  685,  686+2048
,  687,  688,  689,  690+2048
,  691,  692,  693,  694+2048
,  695,  696,  697,  698+2048
,  702,  703,  704,  705+2048
,  706,  707,  708,  709+2048
,  710,  711,  712,  713+2048
,  714,  715,  716,  717+2048
,  718,  719,  720,  721+2048
,  722,  723,  724,  725+2048
,  735,  736,  737,  738+2048
,  739,  740,  741,  742+2048
,  743,  744,  745,  746+2048
,  747,  748,  749,  750+2048
,  754,  755,  756,  757+2048
,  758,  759,  760,  761+2048
,  762,  763,  764,  765+2048
,  766,  767,  768,  769+2048
,  770,  771,  772,  773+2048
,  783,  784,  785,  786+2048
,  790,  791,  792,  793+2048
,  794,  795,  796,  797+2048
,  798,  799,  800,  801+2048
,  802,  803,  804,  805+2048
,  806,  807,  808,  809+2048
,  810,  811,  812,  813+2048
,  814,  815,  816,  817+2048
,  818,  819,  820,  821+2048
,  822,  823,  824,  825+2048
,  826,  827,  828,  829+2048
,  830,  831,  832,  833+2048
,  837,  838,  839,  840+2048
,  841,  842,  843,  844+2048
,  845,  846,  847,  848+2048
,  849,  850,  851,  852+2048
,  853,  854,  855,  856+2048
,  857,  858,  859,  860+2048
,  870,  871,  872,  873+2048
,  874,  875,  876,  877+2048
,  878,  879,  880,  881+2048
,  882,  883,  884,  885+2048
,  889,  890,  891,  892+2048
,  893,  894,  895,  896+2048
,  897,  898,  899,  900+2048
,  901,  902,  903,  904+2048
,  905,  906,  907,  908+2048
,  918,  919,  920,  921+2048
,  925,  926,  927,  928+2048
,  929,  930,  931,  932+2048
,  933,  934,  935,  936+2048
,  937,  938,  939,  940+2048
,  941,  942,  943,  944+2048
,  945,  946,  947,  948+2048
,  949,  950,  951,  952+2048
,  953,  954,  955,  956+2048
,  957,  958,  959,  960+2048
,  961,  962,  963,  964+2048
,  965,  966,  967,  968+2048
,  972,  973,  974,  975+2048
,  976,  977,  978,  979+2048
,  980,  981,  982,  983+2048
,  984,  985,  986,  987+2048
,  988,  989,  990,  991+2048
,  992,  993,  994,  995+2048
, 1005, 1006, 1007, 1008+2048
, 1009, 1010, 1011, 1012+2048
, 1013, 1014, 1015, 1016+2048
, 1017, 1018, 1019, 1020+2048
, 1024, 1025, 1026, 1027+2048
, 1028, 1029, 1030, 1031+2048
, 1032, 1033, 1034, 1035+2048
, 1036, 1037, 1038, 1039+2048
, 1040, 1041, 1042, 1043+2048
, 1053, 1054, 1055, 1056+2048
, 1060, 1061, 1062, 1063+2048
, 1064, 1065, 1066, 1067+2048
, 1068, 1069, 1070, 1071+2048
, 1072, 1073, 1074, 1075+2048
, 1076, 1077, 1078, 1079+2048

,    0,    1,    2,    3,    4+2048
,    5,    6,    7,    8,    9+2048
,   10,   11,   12,   13,   14+2048
,   15,   16,   17,   18,   19+2048
,   20,   21,   22,   23,   24+2048
,   25,   26,   27,   28,   29+2048
,   30,   31,   32,   33,   34+2048
,   35,   36,   37,   38,   39+2048
,   40,   41,   42,   43,   44+2048
,   45,   46,   47,   48,   49+2048
,   50,   51,   52,   53,   54+2048
,   55,   56,   57,   58,   59+2048
,   60,   61,   62,   63,   64+2048
,   65,   66,   67,   68,   69+2048
,   70,   71,   72,   73,   74+2048
,   75,   76,   77,   78,   79+2048
,   80,   81,   82,   83,   84+2048
,   85,   86,   87,   88,   89+2048
,   90,   91,   92,   93,   94+2048
,   95,   96,   97,   98,   99+2048
,  100,  101,  102,  103,  104+2048
,  105,  106,  107,  108,  109+2048
,  110,  111,  112,  113,  114+2048
,  115,  116,  117,  118,  119+2048
,  120,  121,  122,  123,  124+2048
,  125,  126,  127,  128,  129+2048
,  130,  131,  132,  133,  134+2048
,  135,  136,  137,  138,  139+2048
,  140,  141,  142,  143,  144+2048
,  145,  146,  147,  148,  149+2048
,  150,  151,  152,  153,  154+2048
,  155,  156,  157,  158,  159+2048
,  160,  161,  162,  163,  164+2048
,  165,  166,  167,  168,  169+2048
,  170,  171,  172,  173,  174+2048
,  175,  176,  177,  178,  179+2048
,  180,  181,  182,  183,  184+2048
,  185,  186,  187,  188,  189+2048
,  190,  191,  192,  193,  194+2048
,  195,  196,  197,  198,  199+2048
,  200,  201,  202,  203,  204+2048
,  205,  206,  207,  208,  209+2048
,  210,  211,  212,  213,  214+2048
,  215,  216,  217,  218,  219+2048
,  220,  221,  222,  223,  224+2048
,  225,  226,  227,  228,  229+2048
,  230,  231,  232,  233,  234+2048
,  235,  236,  237,  238,  239+2048
,  240,  241,  242,  243,  244+2048
,  245,  246,  247,  248,  249+2048
,  250,  251,  252,  253,  254+2048
,  255,  256,  257,  258,  259+2048
,  260,  261,  262,  263,  264+2048
,  265,  266,  267,  268,  269+2048
,  270,  271,  272,  273,  274+2048
,  275,  276,  277,  278,  279+2048
,  280,  281,  282,  283,  284+2048
,  285,  286,  287,  288,  289+2048
,  290,  291,  292,  293,  294+2048
,  295,  296,  297,  298,  299+2048
,  300,  301,  302,  303,  304+2048
,  305,  306,  307,  308,  309+2048
,  310,  311,  312,  313,  314+2048
,  315,  316,  317,  318,  319+2048
,  320,  321,  322,  323,  324+2048
,  325,  326,  327,  328,  329+2048
,  330,  331,  332,  333,  334+2048
,  335,  336,  337,  338,  339+2048
,  340,  341,  342,  343,  344+2048
,  345,  346,  347,  348,  349+2048
,  350,  351,  352,  353,  354+2048
,  355,  356,  357,  358,  359+2048
,  360,  361,  362,  363,  364+2048
,  365,  366,  367,  368,  369+2048
,  370,  371,  372,  373,  374+2048
,  375,  376,  377,  378,  379+2048
,  380,  381,  382,  383,  384+2048
,  385,  386,  387,  388,  389+2048
,  390,  391,  392,  393,  394+2048
,  395,  396,  397,  398,  399+2048
,  400,  401,  402,  403,  404+2048
,  405,  406,  407,  408,  409+2048
,  410,  411,  412,  413,  414+2048
,  415,  416,  417,  418,  419+2048
,  420,  421,  422,  423,  424+2048
,  425,  426,  427,  428,  429+2048
,  430,  431,  432,  433,  434+2048
,  435,  436,  437,  438,  439+2048
,  440,  441,  442,  443,  444+2048
,  445,  446,  447,  448,  449+2048
,  450,  451,  452,  453,  454+2048
,  455,  456,  457,  458,  459+2048
,  460,  461,  462,  463,  464+2048
,  465,  466,  467,  468,  469+2048
,  470,  471,  472,  473,  474+2048
,  475,  476,  477,  478,  479+2048
,  480,  481,  482,  483,  484+2048
,  485,  486,  487,  488,  489+2048
,  490,  491,  492,  493,  494+2048
,  495,  496,  497,  498,  499+2048
,  500,  501,  502,  503,  504+2048
,  505,  506,  507,  508,  509+2048
,  510,  511,  512,  513,  514+2048
,  515,  516,  517,  518,  519+2048
,  520,  521,  522,  523,  524+2048
,  525,  526,  527,  528,  529+2048
,  530,  531,  532,  533,  534+2048
,  535,  536,  537,  538,  539+2048
,  540,  541,  542,  543,  544+2048
,  545,  546,  547,  548,  549+2048
,  550,  551,  552,  553,  554+2048
,  555,  556,  557,  558,  559+2048
,  560,  561,  562,  563,  564+2048
,  565,  566,  567,  568,  569+2048
,  570,  571,  572,  573,  574+2048
,  575,  576,  577,  578,  579+2048
,  580,  581,  582,  583,  584+2048
,  585,  586,  587,  588,  589+2048
,  590,  591,  592,  593,  594+2048
,  595,  596,  597,  598,  599+2048
,  600,  601,  602,  603,  604+2048
,  605,  606,  607,  608,  609+2048
,  610,  611,  612,  613,  614+2048
,  615,  616,  617,  618,  619+2048
,  620,  621,  622,  623,  624+2048
,  625,  626,  627,  628,  629+2048
,  630,  631,  632,  633,  634+2048
,  635,  636,  637,  638,  639+2048
,  640,  641,  642,  643,  644+2048
,  645,  646,  647,  648,  649+2048
,  650,  651,  652,  653,  654+2048
,  655,  656,  657,  658,  659+2048
,  660,  661,  662,  663,  664+2048
,  665,  666,  667,  668,  669+2048
,  670,  671,  672,  673,  674+2048
,  675,  676,  677,  678,  679+2048
,  680,  681,  682,  683,  684+2048
,  685,  686,  687,  688,  689+2048
,  690,  691,  692,  693,  694+2048
,  695,  696,  697,  698,  699+2048
,  700,  701,  702,  703,  704+2048
,  705,  706,  707,  708,  709+2048
,  710,  711,  712,  713,  714+2048
,  715,  716,  717,  718,  719+2048
,  720,  721,  722,  723,  724+2048
,  725,  726,  727,  728,  729+2048
,  730,  731,  732,  733,  734+2048
,  735,  736,  737,  738,  739+2048
,  740,  741,  742,  743,  744+2048
,  745,  746,  747,  748,  749+2048
,  750,  751,  752,  753,  754+2048
,  755,  756,  757,  758,  759+2048
,  760,  761,  762,  763,  764+2048
,  765,  766,  767,  768,  769+2048
,  770,  771,  772,  773,  774+2048
,  775,  776,  777,  778,  779+2048
,  780,  781,  782,  783,  784+2048
,  785,  786,  787,  788,  789+2048
,  790,  791,  792,  793,  794+2048
,  795,  796,  797,  798,  799+2048
,  800,  801,  802,  803,  804+2048
,  805,  806,  807,  808,  809+2048
,  810,  811,  812,  813,  814+2048
,  815,  816,  817,  818,  819+2048
,  820,  821,  822,  823,  824+2048
,  825,  826,  827,  828,  829+2048
,  830,  831,  832,  833,  834+2048
,  835,  836,  837,  838,  839+2048
,  840,  841,  842,  843,  844+2048
,  845,  846,  847,  848,  849+2048
,  850,  851,  852,  853,  854+2048
,  855,  856,  857,  858,  859+2048
,  860,  861,  862,  863,  864+2048
,  865,  866,  867,  868,  869+2048
,  870,  871,  872,  873,  874+2048
,  875,  876,  877,  878,  879+2048
,  880,  881,  882,  883,  884+2048
,  885,  886,  887,  888,  889+2048
,  890,  891,  892,  893,  894+2048
,  895,  896,  897,  898,  899+2048
,  900,  901,  902,  903,  904+2048
,  905,  906,  907,  908,  909+2048
,  910,  911,  912,  913,  914+2048
,  915,  916,  917,  918,  919+2048
,  920,  921,  922,  923,  924+2048
,  925,  926,  927,  928,  929+2048
,  930,  931,  932,  933,  934+2048
,  935,  936,  937,  938,  939+2048
,  940,  941,  942,  943,  944+2048
,  945,  946,  947,  948,  949+2048
,  950,  951,  952,  953,  954+2048
,  955,  956,  957,  958,  959+2048
,  960,  961,  962,  963,  964+2048
,  965,  966,  967,  968,  969+2048
,  970,  971,  972,  973,  974+2048
,  975,  976,  977,  978,  979+2048
,  980,  981,  982,  983,  984+2048
,  985,  986,  987,  988,  989+2048
,  990,  991,  992,  993,  994+2048
,  995,  996,  997,  998,  999+2048
, 1000, 1001, 1002, 1003, 1004+2048
, 1005, 1006, 1007, 1008, 1009+2048
, 1010, 1011, 1012, 1013, 1014+2048
, 1015, 1016, 1017, 1018, 1019+2048
, 1020, 1021, 1022, 1023, 1024+2048
, 1025, 1026, 1027, 1028, 1029+2048
, 1030, 1031, 1032, 1033, 1034+2048
, 1035, 1036, 1037, 1038, 1039+2048
, 1040, 1041, 1042, 1043, 1044+2048
, 1045, 1046, 1047, 1048, 1049+2048
, 1050, 1051, 1052, 1053, 1054+2048
, 1055, 1056, 1057, 1058, 1059+2048
, 1060, 1061, 1062, 1063, 1064+2048
, 1065, 1066, 1067, 1068, 1069+2048
, 1070, 1071, 1072, 1073, 1074+2048
, 1075, 1076, 1077, 1078, 1079+2048
, 1080, 1081, 1082, 1083, 1084+2048
, 1085, 1086, 1087, 1088, 1089+2048
, 1090, 1091, 1092, 1093, 1094+2048
, 1095, 1096, 1097, 1098, 1099+2048
, 1100, 1101, 1102, 1103, 1104+2048
, 1105, 1106, 1107, 1108, 1109+2048
, 1110, 1111, 1112, 1113, 1114+2048
, 1115, 1116, 1117, 1118, 1119+2048
, 1120, 1121, 1122, 1123, 1124+2048
, 1125, 1126, 1127, 1128, 1129+2048
, 1130, 1131, 1132, 1133, 1134+2048
, 1135, 1136, 1137, 1138, 1139+2048
, 1140, 1141, 1142, 1143, 1144+2048
, 1145, 1146, 1147, 1148, 1149+2048
, 1150, 1151, 1152, 1153, 1154+2048
, 1155, 1156, 1157, 1158, 1159+2048
, 1160, 1161, 1162, 1163, 1164+2048
, 1165, 1166, 1167, 1168, 1169+2048
, 1170, 1171, 1172, 1173, 1174+2048
, 1175, 1176, 1177, 1178, 1179+2048
, 1180, 1181, 1182, 1183, 1184+2048
, 1185, 1186, 1187, 1188, 1189+2048
, 1190, 1191, 1192, 1193, 1194+2048
, 1195, 1196, 1197, 1198, 1199+2048

,    0,    1,    2,    3,    4,    5+2048
,    6,    7,    8,    9,   10,   11+2048
,   12,   13,   14,   15,   16,   17+2048
,   18,   19,   20,   21,   22,   23+2048
,   24,   25,   26,   27,   28,   29+2048
,   30,   31,   32,   33,   34,   35+2048
,   36,   37,   38,   39,   40,   41+2048
,   42,   43,   44,   45,   46,   47+2048
,   48,   49,   50,   51,   52,   53+2048
,   54,   55,   56,   57,   58,   59+2048
,   60,   61,   62,   63,   64,   65+2048
,   66,   67,   68,   69,   70,   71+2048
,   72,   73,   74,   75,   76,   77+2048
,   78,   79,   80,   81,   82,   83+2048
,   84,   85,   86,   87,   88,   89+2048
,   90,   91,   92,   93,   94,   95+2048
,   96,   97,   98,   99,  100,  101+2048
,  102,  103,  104,  105,  106,  107+2048
,  108,  109,  110,  111,  112,  113+2048
,  114,  115,  116,  117,  118,  119+2048
,  120,  121,  122,  123,  124,  125+2048
,  126,  127,  128,  129,  130,  131+2048
,  132,  133,  134,  135,  136,  137+2048
,  138,  139,  140,  141,  142,  143+2048
,  144,  145,  146,  147,  148,  149+2048
,  150,  151,  152,  153,  154,  155+2048
,  156,  157,  158,  159,  160,  161+2048
,  162,  163,  164,  165,  166,  167+2048
,  168,  169,  170,  171,  172,  173+2048
,  174,  175,  176,  177,  178,  179+2048
,  180,  181,  182,  183,  184,  185+2048
,  186,  187,  188,  189,  190,  191+2048
,  192,  193,  194,  195,  196,  197+2048
,  198,  199,  200,  201,  202,  203+2048
,  204,  205,  206,  207,  208,  209+2048
,  210,  211,  212,  213,  214,  215+2048
,  216,  217,  218,  219,  220,  221+2048
,  222,  223,  224,  225,  226,  227+2048
,  228,  229,  230,  231,  232,  233+2048
,  234,  235,  236,  237,  238,  239+2048
,  240,  241,  242,  243,  244,  245+2048
,  246,  247,  248,  249,  250,  251+2048
,  252,  253,  254,  255,  256,  257+2048
,  258,  259,  260,  261,  262,  263+2048
,  264,  265,  266,  267,  268,  269+2048
,  270,  271,  272,  273,  274,  275+2048
,  276,  277,  278,  279,  280,  281+2048
,  282,  283,  284,  285,  286,  287+2048
,  288,  289,  290,  291,  292,  293+2048
,  294,  295,  296,  297,  298,  299+2048
,  300,  301,  302,  303,  304,  305+2048
,  306,  307,  308,  309,  310,  311+2048
,  312,  313,  314,  315,  316,  317+2048
,  318,  319,  320,  321,  322,  323+2048
,  324,  325,  326,  327,  328,  329+2048
,  330,  331,  332,  333,  334,  335+2048
,  336,  337,  338,  339,  340,  341+2048
,  342,  343,  344,  345,  346,  347+2048
,  348,  349,  350,  351,  352,  353+2048
,  354,  355,  356,  357,  358,  359+2048
,  360,  361,  362,  363,  364,  365+2048
,  366,  367,  368,  369,  370,  371+2048
,  372,  373,  374,  375,  376,  377+2048
,  378,  379,  380,  381,  382,  383+2048
,  384,  385,  386,  387,  388,  389+2048
,  390,  391,  392,  393,  394,  395+2048
,  396,  397,  398,  399,  400,  401+2048
,  402,  403,  404,  405,  406,  407+2048
,  408,  409,  410,  411,  412,  413+2048
,  414,  415,  416,  417,  418,  419+2048
,  420,  421,  422,  423,  424,  425+2048
,  426,  427,  428,  429,  430,  431+2048
,  432,  433,  434,  435,  436,  437+2048
,  438,  439,  440,  441,  442,  443+2048
,  444,  445,  446,  447,  448,  449+2048
,  450,  451,  452,  453,  454,  455+2048
,  456,  457,  458,  459,  460,  461+2048
,  462,  463,  464,  465,  466,  467+2048
,  468,  469,  470,  471,  472,  473+2048
,  474,  475,  476,  477,  478,  479+2048
,  480,  481,  482,  483,  484,  485+2048
,  486,  487,  488,  489,  490,  491+2048
,  492,  493,  494,  495,  496,  497+2048
,  498,  499,  500,  501,  502,  503+2048
,  504,  505,  506,  507,  508,  509+2048
,  510,  511,  512,  513,  514,  515+2048
,  516,  517,  518,  519,  520,  521+2048
,  522,  523,  524,  525,  526,  527+2048
,  528,  529,  530,  531,  532,  533+2048
,  534,  535,  536,  537,  538,  539+2048
,  540,  541,  542,  543,  544,  545+2048
,  546,  547,  548,  549,  550,  551+2048
,  552,  553,  554,  555,  556,  557+2048
,  558,  559,  560,  561,  562,  563+2048
,  564,  565,  566,  567,  568,  569+2048
,  570,  571,  572,  573,  574,  575+2048
,  576,  577,  578,  579,  580,  581+2048
,  582,  583,  584,  585,  586,  587+2048
,  588,  589,  590,  591,  592,  593+2048
,  594,  595,  596,  597,  598,  599+2048
,  600,  601,  602,  603,  604,  605+2048
,  606,  607,  608,  609,  610,  611+2048
,  612,  613,  614,  615,  616,  617+2048
,  618,  619,  620,  621,  622,  623+2048
,  624,  625,  626,  627,  628,  629+2048
,  630,  631,  632,  633,  634,  635+2048
,  636,  637,  638,  639,  640,  641+2048
,  642,  643,  644,  645,  646,  647+2048
,  648,  649,  650,  651,  652,  653+2048
,  654,  655,  656,  657,  658,  659+2048
,  660,  661,  662,  663,  664,  665+2048
,  666,  667,  668,  669,  670,  671+2048
,  672,  673,  674,  675,  676,  677+2048
,  678,  679,  680,  681,  682,  683+2048
,  684,  685,  686,  687,  688,  689+2048
,  690,  691,  692,  693,  694,  695+2048
,  696,  697,  698,  699,  700,  701+2048
,  702,  703,  704,  705,  706,  707+2048
,  708,  709,  710,  711,  712,  713+2048
,  714,  715,  716,  717,  718,  719+2048
,  720,  721,  722,  723,  724,  725+2048
,  726,  727,  728,  729,  730,  731+2048
,  732,  733,  734,  735,  736,  737+2048
,  738,  739,  740,  741,  742,  743+2048
,  744,  745,  746,  747,  748,  749+2048
,  750,  751,  752,  753,  754,  755+2048
,  756,  757,  758,  759,  760,  761+2048
,  762,  763,  764,  765,  766,  767+2048
,  768,  769,  770,  771,  772,  773+2048
,  774,  775,  776,  777,  778,  779+2048
,  780,  781,  782,  783,  784,  785+2048
,  786,  787,  788,  789,  790,  791+2048
,  792,  793,  794,  795,  796,  797+2048
,  798,  799,  800,  801,  802,  803+2048
,  804,  805,  806,  807,  808,  809+2048
,  810,  811,  812,  813,  814,  815+2048
,  816,  817,  818,  819,  820,  821+2048
,  822,  823,  824,  825,  826,  827+2048
,  828,  829,  830,  831,  832,  833+2048
,  834,  835,  836,  837,  838,  839+2048
,  840,  841,  842,  843,  844,  845+2048
,  846,  847,  848,  849,  850,  851+2048
,  852,  853,  854,  855,  856,  857+2048
,  858,  859,  860,  861,  862,  863+2048
,  864,  865,  866,  867,  868,  869+2048
,  870,  871,  872,  873,  874,  875+2048
,  876,  877,  878,  879,  880,  881+2048
,  882,  883,  884,  885,  886,  887+2048
,  888,  889,  890,  891,  892,  893+2048
,  894,  895,  896,  897,  898,  899+2048
,  900,  901,  902,  903,  904,  905+2048
,  906,  907,  908,  909,  910,  911+2048
,  912,  913,  914,  915,  916,  917+2048
,  918,  919,  920,  921,  922,  923+2048
,  924,  925,  926,  927,  928,  929+2048
,  930,  931,  932,  933,  934,  935+2048
,  936,  937,  938,  939,  940,  941+2048
,  942,  943,  944,  945,  946,  947+2048
,  948,  949,  950,  951,  952,  953+2048
,  954,  955,  956,  957,  958,  959+2048
,  960,  961,  962,  963,  964,  965+2048
,  966,  967,  968,  969,  970,  971+2048
,  972,  973,  974,  975,  976,  977+2048
,  978,  979,  980,  981,  982,  983+2048
,  984,  985,  986,  987,  988,  989+2048
,  990,  991,  992,  993,  994,  995+2048
,  996,  997,  998,  999, 1000, 1001+2048
, 1002, 1003, 1004, 1005, 1006, 1007+2048
, 1008, 1009, 1010, 1011, 1012, 1013+2048
, 1014, 1015, 1016, 1017, 1018, 1019+2048
, 1020, 1021, 1022, 1023, 1024, 1025+2048
, 1026, 1027, 1028, 1029, 1030, 1031+2048
, 1032, 1033, 1034, 1035, 1036, 1037+2048
, 1038, 1039, 1040, 1041, 1042, 1043+2048
, 1044, 1045, 1046, 1047, 1048, 1049+2048
, 1050, 1051, 1052, 1053, 1054, 1055+2048
, 1056, 1057, 1058, 1059, 1060, 1061+2048
, 1062, 1063, 1064, 1065, 1066, 1067+2048
, 1068, 1069, 1070, 1071, 1072, 1073+2048
, 1074, 1075, 1076, 1077, 1078, 1079+2048
, 1080, 1081, 1082, 1083, 1084, 1085+2048
, 1086, 1087, 1088, 1089, 1090, 1091+2048
, 1092, 1093, 1094, 1095, 1096, 1097+2048
, 1098, 1099, 1100, 1101, 1102, 1103+2048
, 1104, 1105, 1106, 1107, 1108, 1109+2048
, 1110, 1111, 1112, 1113, 1114, 1115+2048
, 1116, 1117, 1118, 1119, 1120, 1121+2048
, 1122, 1123, 1124, 1125, 1126, 1127+2048
, 1128, 1129, 1130, 1131, 1132, 1133+2048
, 1134, 1135, 1136, 1137, 1138, 1139+2048
, 1140, 1141, 1142, 1143, 1144, 1145+2048
, 1146, 1147, 1148, 1149, 1150, 1151+2048
, 1152, 1153, 1154, 1155, 1156, 1157+2048
, 1158, 1159, 1160, 1161, 1162, 1163+2048
, 1164, 1165, 1166, 1167, 1168, 1169+2048
, 1170, 1171, 1172, 1173, 1174, 1175+2048
, 1176, 1177, 1178, 1179, 1180, 1181+2048
, 1182, 1183, 1184, 1185, 1186, 1187+2048
, 1188, 1189, 1190, 1191, 1192, 1193+2048
, 1194, 1195, 1196, 1197, 1198, 1199+2048
, 1200, 1201, 1202, 1203, 1204, 1205+2048
, 1206, 1207, 1208, 1209, 1210, 1211+2048
, 1212, 1213, 1214, 1215, 1216, 1217+2048
, 1218, 1219, 1220, 1221, 1222, 1223+2048
, 1224, 1225, 1226, 1227, 1228, 1229+2048
, 1230, 1231, 1232, 1233, 1234, 1235+2048
, 1236, 1237, 1238, 1239, 1240, 1241+2048
, 1242, 1243, 1244, 1245, 1246, 1247+2048
, 1248, 1249, 1250, 1251, 1252, 1253+2048
, 1254, 1255, 1256, 1257, 1258, 1259+2048
, 1260, 1261, 1262, 1263, 1264, 1265+2048
, 1266, 1267, 1268, 1269, 1270, 1271+2048
, 1272, 1273, 1274, 1275, 1276, 1277+2048
, 1278, 1279, 1280, 1281, 1282, 1283+2048
, 1284, 1285, 1286, 1287, 1288, 1289+2048
, 1290, 1291, 1292, 1293, 1294, 1295+2048

,   24,   25,   26,   27+2048
,   33,   34,   35,   36+2048
,   87,   88,   89,   90+2048
,  102,  103,  104,  105+2048
,  159,  160,  161,  162+2048
,  168,  169,  170,  171+2048
,  222,  223,  224,  225+2048
,  237,  238,  239,  240+2048
,  294,  295,  296,  297+2048
,  303,  304,  305,  306+2048
,  357,  358,  359,  360+2048
,  372,  373,  374,  375+2048
,  429,  430,  431,  432+2048
,  438,  439,  440,  441+2048
,  492,  493,  494,  495+2048
,  507,  508,  509,  510+2048
,  564,  565,  566,  567+2048
,  573,  574,  575,  576+2048
,  627,  628,  629,  630+2048
,  642,  643,  644,  645+2048
,  699,  700,  701,  702+2048
,  708,  709,  710,  711+2048
,  762,  763,  764,  765+2048
,  777,  778,  779,  780+2048
,  834,  835,  836,  837+2048
,  843,  844,  845,  846+2048
,  897,  898,  899,  900+2048
,  912,  913,  914,  915+2048
,  969,  970,  971,  972+2048
,  978,  979,  980,  981+2048
, 1032, 1033, 1034, 1035+2048
, 1047, 1048, 1049, 1050+2048
,    0,    1,    2,    3,    4+2048
,   28,   29,   30,   31,   32+2048
,   37,   38,   39,   40,   41+2048
,   48,   49,   50,   51,   52+2048
,   53,   54,   55,   56,   57+2048
,   82,   83,   84,   85,   86+2048
,   97,   98,   99,  100,  101+2048
,  112,  113,  114,  115,  116+2048
,  123,  124,  125,  126,  127+2048
,  135,  136,  137,  138,  139+2048
,  163,  164,  165,  166,  167+2048
,  172,  173,  174,  175,  176+2048
,  183,  184,  185,  186,  187+2048
,  188,  189,  190,  191,  192+2048
,  217,  218,  219,  220,  221+2048
,  232,  233,  234,  235,  236+2048
,  247,  248,  249,  250,  251+2048
,  258,  259,  260,  261,  262+2048
,  270,  271,  272,  273,  274+2048
,  298,  299,  300,  301,  302+2048
,  307,  308,  309,  310,  311+2048
,  318,  319,  320,  321,  322+2048
,  323,  324,  325,  326,  327+2048
,  352,  353,  354,  355,  356+2048
,  367,  368,  369,  370,  371+2048
,  382,  383,  384,  385,  386+2048
,  393,  394,  395,  396,  397+2048
,  405,  406,  407,  408,  409+2048
,  433,  434,  435,  436,  437+2048
,  442,  443,  444,  445,  446+2048
,  453,  454,  455,  456,  457+2048
,  458,  459,  460,  461,  462+2048
,  487,  488,  489,  490,  491+2048
,  502,  503,  504,  505,  506+2048
,  517,  518,  519,  520,  521+2048
,  528,  529,  530,  531,  532+2048
,  540,  541,  542,  543,  544+2048
,  568,  569,  570,  571,  572+2048
,  577,  578,  579,  580,  581+2048
,  588,  589,  590,  591,  592+2048
,  593,  594,  595,  596,  597+2048
,  622,  623,  624,  625,  626+2048
,  637,  638,  639,  640,  641+2048
,  652,  653,  654,  655,  656+2048
,  663,  664,  665,  666,  667+2048
,  675,  676,  677,  678,  679+2048
,  703,  704,  705,  706,  707+2048
,  712,  713,  714,  715,  716+2048
,  723,  724,  725,  726,  727+2048
,  728,  729,  730,  731,  732+2048
,  757,  758,  759,  760,  761+2048
,  772,  773,  774,  775,  776+2048
,  787,  788,  789,  790,  791+2048
,  798,  799,  800,  801,  802+2048
,  810,  811,  812,  813,  814+2048
,  838,  839,  840,  841,  842+2048
,  847,  848,  849,  850,  851+2048
,  858,  859,  860,  861,  862+2048
,  863,  864,  865,  866,  867+2048
,  892,  893,  894,  895,  896+2048
,  907,  908,  909,  910,  911+2048
,  922,  923,  924,  925,  926+2048
,  933,  934,  935,  936,  937+2048
,  945,  946,  947,  948,  949+2048
,  973,  974,  975,  976,  977+2048
,  982,  983,  984,  985,  986+2048
,  993,  994,  995,  996,  997+2048
,  998,  999, 1000, 1001, 1002+2048
, 1027, 1028, 1029, 1030, 1031+2048
, 1042, 1043, 1044, 1045, 1046+2048
, 1057, 1058, 1059, 1060, 1061+2048
, 1068, 1069, 1070, 1071, 1072+2048
,    5,    6,    7,    8,    9,   10+2048
,   18,   19,   20,   21,   22,   23+2048
,   42,   43,   44,   45,   46,   47+2048
,   58,   59,   60,   61,   62,   63+2048
,   64,   65,   66,   67,   68,   69+2048
,   70,   71,   72,   73,   74,   75+2048
,   76,   77,   78,   79,   80,   81+2048
,   91,   92,   93,   94,   95,   96+2048
,  106,  107,  108,  109,  110,  111+2048
,  117,  118,  119,  120,  121,  122+2048
,  140,  141,  142,  143,  144,  145+2048
,  153,  154,  155,  156,  157,  158+2048
,  177,  178,  179,  180,  181,  182+2048
,  193,  194,  195,  196,  197,  198+2048
,  199,  200,  201,  202,  203,  204+2048
,  205,  206,  207,  208,  209,  210+2048
,  211,  212,  213,  214,  215,  216+2048
,  226,  227,  228,  229,  230,  231+2048
,  241,  242,  243,  244,  245,  246+2048
,  252,  253,  254,  255,  256,  257+2048
,  275,  276,  277,  278,  279,  280+2048
,  288,  289,  290,  291,  292,  293+2048
,  312,  313,  314,  315,  316,  317+2048
,  328,  329,  330,  331,  332,  333+2048
,  334,  335,  336,  337,  338,  339+2048
,  340,  341,  342,  343,  344,  345+2048
,  346,  347,  348,  349,  350,  351+2048
,  361,  362,  363,  364,  365,  366+2048
,  376,  377,  378,  379,  380,  381+2048
,  387,  388,  389,  390,  391,  392+2048
,  410,  411,  412,  413,  414,  415+2048
,  423,  424,  425,  426,  427,  428+2048
,  447,  448,  449,  450,  451,  452+2048
,  463,  464,  465,  466,  467,  468+2048
,  469,  470,  471,  472,  473,  474+2048
,  475,  476,  477,  478,  479,  480+2048
,  481,  482,  483,  484,  485,  486+2048
,  496,  497,  498,  499,  500,  501+2048
,  511,  512,  513,  514,  515,  516+2048
,  522,  523,  524,  525,  526,  527+2048
,  545,  546,  547,  548,  549,  550+2048
,  558,  559,  560,  561,  562,  563+2048
,  582,  583,  584,  585,  586,  587+2048
,  598,  599,  600,  601,  602,  603+2048
,  604,  605,  606,  607,  608,  609+2048
,  610,  611,  612,  613,  614,  615+2048
,  616,  617,  618,  619,  620,  621+2048
,  631,  632,  633,  634,  635,  636+2048
,  646,  647,  648,  649,  650,  651+2048
,  657,  658,  659,  660,  661,  662+2048
,  680,  681,  682,  683,  684,  685+2048
,  693,  694,  695,  696,  697,  698+2048
,  717,  718,  719,  720,  721,  722+2048
,  733,  734,  735,  736,  737,  738+2048
,  739,  740,  741,  742,  743,  744+2048
,  745,  746,  747,  748,  749,  750+2048
,  751,  752,  753,  754,  755,  756+2048
,  766,  767,  768,  769,  770,  771+2048
,  781,  782,  783,  784,  785,  786+2048
,  792,  793,  794,  795,  796,  797+2048
,  815,  816,  817,  818,  819,  820+2048
,  828,  829,  830,  831,  832,  833+2048
,  852,  853,  854,  855,  856,  857+2048
,  868,  869,  870,  871,  872,  873+2048
,  874,  875,  876,  877,  878,  879+2048
,  880,  881,  882,  883,  884,  885+2048
,  886,  887,  888,  889,  890,  891+2048
,  901,  902,  903,  904,  905,  906+2048
,  916,  917,  918,  919,  920,  921+2048
,  927,  928,  929,  930,  931,  932+2048
,  950,  951,  952,  953,  954,  955+2048
,  963,  964,  965,  966,  967,  968+2048
,  987,  988,  989,  990,  991,  992+2048
, 1003, 1004, 1005, 1006, 1007, 1008+2048
, 1009, 1010, 1011, 1012, 1013, 1014+2048
, 1015, 1016, 1017, 1018, 1019, 1020+2048
, 1021, 1022, 1023, 1024, 1025, 1026+2048
, 1036, 1037, 1038, 1039, 1040, 1041+2048
, 1051, 1052, 1053, 1054, 1055, 1056+2048
, 1062, 1063, 1064, 1065, 1066, 1067+2048
,   11,   12,   13,   14,   15,   16,   17+2048
,  128,  129,  130,  131,  132,  133,  134+2048
,  146,  147,  148,  149,  150,  151,  152+2048
,  263,  264,  265,  266,  267,  268,  269+2048
,  281,  282,  283,  284,  285,  286,  287+2048
,  398,  399,  400,  401,  402,  403,  404+2048
,  416,  417,  418,  419,  420,  421,  422+2048
,  533,  534,  535,  536,  537,  538,  539+2048
,  551,  552,  553,  554,  555,  556,  557+2048
,  668,  669,  670,  671,  672,  673,  674+2048
,  686,  687,  688,  689,  690,  691,  692+2048
,  803,  804,  805,  806,  807,  808,  809+2048
,  821,  822,  823,  824,  825,  826,  827+2048
,  938,  939,  940,  941,  942,  943,  944+2048
,  956,  957,  958,  959,  960,  961,  962+2048
, 1073, 1074, 1075, 1076, 1077, 1078, 1079+2048

,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9,   10+2048
,   11,   12,   13,   14,   15,   16,   17,   18,   19,   20,   21+2048
,   22,   23,   24,   25,   26,   27,   28,   29,   30,   31,   32+2048
,   33,   34,   35,   36,   37,   38,   39,   40,   41,   42,   43+2048
,   44,   45,   46,   47,   48,   49,   50,   51,   52,   53,   54+2048
,   55,   56,   57,   58,   59,   60,   61,   62,   63,   64,   65+2048
,   66,   67,   68,   69,   70,   71,   72,   73,   74,   75,   76+2048
,   77,   78,   79,   80,   81,   82,   83,   84,   85,   86,   87+2048
,   88,   89,   90,   91,   92,   93,   94,   95,   96,   97,   98+2048
,   99,  100,  101,  102,  103,  104,  105,  106,  107,  108,  109+2048
,  110,  111,  112,  113,  114,  115,  116,  117,  118,  119,  120+2048
,  121,  122,  123,  124,  125,  126,  127,  128,  129,  130,  131+2048
,  132,  133,  134,  135,  136,  137,  138,  139,  140,  141,  142+2048
,  143,  144,  145,  146,  147,  148,  149,  150,  151,  152,  153+2048
,  154,  155,  156,  157,  158,  159,  160,  161,  162,  163,  164+2048
,  165,  166,  167,  168,  169,  170,  171,  172,  173,  174,  175+2048
,  176,  177,  178,  179,  180,  181,  182,  183,  184,  185,  186+2048
,  187,  188,  189,  190,  191,  192,  193,  194,  195,  196,  197+2048
,  198,  199,  200,  201,  202,  203,  204,  205,  206,  207,  208+2048
,  209,  210,  211,  212,  213,  214,  215,  216,  217,  218,  219+2048
,  220,  221,  222,  223,  224,  225,  226,  227,  228,  229,  230+2048
,  231,  232,  233,  234,  235,  236,  237,  238,  239,  240,  241+2048
,  242,  243,  244,  245,  246,  247,  248,  249,  250,  251,  252+2048
,  253,  254,  255,  256,  257,  258,  259,  260,  261,  262,  263+2048
,  264,  265,  266,  267,  268,  269,  270,  271,  272,  273,  274+2048
,  275,  276,  277,  278,  279,  280,  281,  282,  283,  284,  285+2048
,  286,  287,  288,  289,  290,  291,  292,  293,  294,  295,  296+2048
,  297,  298,  299,  300,  301,  302,  303,  304,  305,  306,  307+2048
,  308,  309,  310,  311,  312,  313,  314,  315,  316,  317,  318+2048
,  319,  320,  321,  322,  323,  324,  325,  326,  327,  328,  329+2048
,  330,  331,  332,  333,  334,  335,  336,  337,  338,  339,  340+2048
,  341,  342,  343,  344,  345,  346,  347,  348,  349,  350,  351+2048
,  352,  353,  354,  355,  356,  357,  358,  359,  360,  361,  362+2048
,  363,  364,  365,  366,  367,  368,  369,  370,  371,  372,  373+2048
,  374,  375,  376,  377,  378,  379,  380,  381,  382,  383,  384+2048
,  385,  386,  387,  388,  389,  390,  391,  392,  393,  394,  395+2048
,  396,  397,  398,  399,  400,  401,  402,  403,  404,  405,  406+2048
,  407,  408,  409,  410,  411,  412,  413,  414,  415,  416,  417+2048
,  418,  419,  420,  421,  422,  423,  424,  425,  426,  427,  428+2048
,  429,  430,  431,  432,  433,  434,  435,  436,  437,  438,  439+2048
,  440,  441,  442,  443,  444,  445,  446,  447,  448,  449,  450+2048
,  451,  452,  453,  454,  455,  456,  457,  458,  459,  460,  461+2048
,  462,  463,  464,  465,  466,  467,  468,  469,  470,  471,  472+2048
,  473,  474,  475,  476,  477,  478,  479,  480,  481,  482,  483+2048
,  484,  485,  486,  487,  488,  489,  490,  491,  492,  493,  494+2048
,  495,  496,  497,  498,  499,  500,  501,  502,  503,  504,  505+2048
,  506,  507,  508,  509,  510,  511,  512,  513,  514,  515,  516+2048
,  517,  518,  519,  520,  521,  522,  523,  524,  525,  526,  527+2048
,  528,  529,  530,  531,  532,  533,  534,  535,  536,  537,  538+2048
,  539,  540,  541,  542,  543,  544,  545,  546,  547,  548,  549+2048
,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559,  560+2048
,  561,  562,  563,  564,  565,  566,  567,  568,  569,  570,  571+2048
,  572,  573,  574,  575,  576,  577,  578,  579,  580,  581,  582+2048
,  583,  584,  585,  586,  587,  588,  589,  590,  591,  592,  593+2048
,  594,  595,  596,  597,  598,  599,  600,  601,  602,  603,  604+2048
,  605,  606,  607,  608,  609,  610,  611,  612,  613,  614,  615+2048
,  616,  617,  618,  619,  620,  621,  622,  623,  624,  625,  626+2048
,  627,  628,  629,  630,  631,  632,  633,  634,  635,  636,  637+2048
,  638,  639,  640,  641,  642,  643,  644,  645,  646,  647,  648+2048
,  649,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659+2048
,  660,  661,  662,  663,  664,  665,  666,  667,  668,  669,  670+2048
,  671,  672,  673,  674,  675,  676,  677,  678,  679,  680,  681+2048
,  682,  683,  684,  685,  686,  687,  688,  689,  690,  691,  692+2048
,  693,  694,  695,  696,  697,  698,  699,  700,  701,  702,  703+2048
,  704,  705,  706,  707,  708,  709,  710,  711,  712,  713,  714+2048
,  715,  716,  717,  718,  719,  720,  721,  722,  723,  724,  725+2048
,  726,  727,  728,  729,  730,  731,  732,  733,  734,  735,  736+2048
,  737,  738,  739,  740,  741,  742,  743,  744,  745,  746,  747+2048
,  748,  749,  750,  751,  752,  753,  754,  755,  756,  757,  758+2048
,  759,  760,  761,  762,  763,  764,  765,  766,  767,  768,  769+2048
,  770,  771,  772,  773,  774,  775,  776,  777,  778,  779,  780+2048
,  781,  782,  783,  784,  785,  786,  787,  788,  789,  790,  791+2048
,  792,  793,  794,  795,  796,  797,  798,  799,  800,  801,  802+2048
,  803,  804,  805,  806,  807,  808,  809,  810,  811,  812,  813+2048
,  814,  815,  816,  817,  818,  819,  820,  821,  822,  823,  824+2048
,  825,  826,  827,  828,  829,  830,  831,  832,  833,  834,  835+2048
,  836,  837,  838,  839,  840,  841,  842,  843,  844,  845,  846+2048
,  847,  848,  849,  850,  851,  852,  853,  854,  855,  856,  857+2048
,  858,  859,  860,  861,  862,  863,  864,  865,  866,  867,  868+2048
,  869,  870,  871,  872,  873,  874,  875,  876,  877,  878,  879+2048
,  880,  881,  882,  883,  884,  885,  886,  887,  888,  889,  890+2048
,  891,  892,  893,  894,  895,  896,  897,  898,  899,  900,  901+2048
,  902,  903,  904,  905,  906,  907,  908,  909,  910,  911,  912+2048
,  913,  914,  915,  916,  917,  918,  919,  920,  921,  922,  923+2048
,  924,  925,  926,  927,  928,  929,  930,  931,  932,  933,  934+2048
,  935,  936,  937,  938,  939,  940,  941,  942,  943,  944,  945+2048
,  946,  947,  948,  949,  950,  951,  952,  953,  954,  955,  956+2048
,  957,  958,  959,  960,  961,  962,  963,  964,  965,  966,  967+2048
,  968,  969,  970,  971,  972,  973,  974,  975,  976,  977,  978+2048
,  979,  980,  981,  982,  983,  984,  985,  986,  987,  988,  989+2048
,  990,  991,  992,  993,  994,  995,  996,  997,  998,  999, 1000+2048
, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011+2048
, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022+2048
, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033+2048
, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044+2048
, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055+2048
, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066+2048
, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077+2048
, 1078, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088+2048
, 1089, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099+2048
, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109, 1110+2048
, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119, 1120, 1121+2048
, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129, 1130, 1131, 1132+2048
, 1133, 1134, 1135, 1136, 1137, 1138, 1139, 1140, 1141, 1142, 1143+2048
, 1144, 1145, 1146, 1147, 1148, 1149, 1150, 1151, 1152, 1153, 1154+2048
, 1155, 1156, 1157, 1158, 1159, 1160, 1161, 1162, 1163, 1164, 1165+2048
, 1166, 1167, 1168, 1169, 1170, 1171, 1172, 1173, 1174, 1175, 1176+2048
, 1177, 1178, 1179, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187+2048
, 1188, 1189, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198+2048
, 1199, 1200, 1201, 1202, 1203, 1204, 1205, 1206, 1207, 1208, 1209+2048
, 1210, 1211, 1212, 1213, 1214, 1215, 1216, 1217, 1218, 1219, 1220+2048
, 1221, 1222, 1223, 1224, 1225, 1226, 1227, 1228, 1229, 1230, 1231+2048
, 1232, 1233, 1234, 1235, 1236, 1237, 1238, 1239, 1240, 1241, 1242+2048
, 1243, 1244, 1245, 1246, 1247, 1248, 1249, 1250, 1251, 1252, 1253+2048
, 1254, 1255, 1256, 1257, 1258, 1259, 1260, 1261, 1262, 1263, 1264+2048
, 1265, 1266, 1267, 1268, 1269, 1270, 1271, 1272, 1273, 1274, 1275+2048
, 1276, 1277, 1278, 1279, 1280, 1281, 1282, 1283, 1284, 1285, 1286+2048
, 1287, 1288, 1289, 1290, 1291, 1292, 1293, 1294, 1295, 1296, 1297+2048
, 1298, 1299, 1300, 1301, 1302, 1303, 1304, 1305, 1306, 1307, 1308+2048
, 1309, 1310, 1311, 1312, 1313, 1314, 1315, 1316, 1317, 1318, 1319+2048
, 1320, 1321, 1322, 1323, 1324, 1325, 1326, 1327, 1328, 1329, 1330+2048
, 1331, 1332, 1333, 1334, 1335, 1336, 1337, 1338, 1339, 1340, 1341+2048
, 1342, 1343, 1344, 1345, 1346, 1347, 1348, 1349, 1350, 1351, 1352+2048
, 1353, 1354, 1355, 1356, 1357, 1358, 1359, 1360, 1361, 1362, 1363+2048
, 1364, 1365, 1366, 1367, 1368, 1369, 1370, 1371, 1372, 1373, 1374+2048
, 1375, 1376, 1377, 1378, 1379, 1380, 1381, 1382, 1383, 1384, 1385+2048
, 1386, 1387, 1388, 1389, 1390, 1391, 1392, 1393, 1394, 1395, 1396+2048
, 1397, 1398, 1399, 1400, 1401, 1402, 1403, 1404, 1405, 1406, 1407+2048
, 1408, 1409, 1410, 1411, 1412, 1413, 1414, 1415, 1416, 1417, 1418+2048
, 1419, 1420, 1421, 1422, 1423, 1424, 1425, 1426, 1427, 1428, 1429+2048
, 1430, 1431, 1432, 1433, 1434, 1435, 1436, 1437, 1438, 1439, 1440+2048
, 1441, 1442, 1443, 1444, 1445, 1446, 1447, 1448, 1449, 1450, 1451+2048
, 1452, 1453, 1454, 1455, 1456, 1457, 1458, 1459, 1460, 1461, 1462+2048
, 1463, 1464, 1465, 1466, 1467, 1468, 1469, 1470, 1471, 1472, 1473+2048
, 1474, 1475, 1476, 1477, 1478, 1479, 1480, 1481, 1482, 1483, 1484+2048
, 1485, 1486, 1487, 1488, 1489, 1490, 1491, 1492, 1493, 1494, 1495+2048
, 1496, 1497, 1498, 1499, 1500, 1501, 1502, 1503, 1504, 1505, 1506+2048
, 1507, 1508, 1509, 1510, 1511, 1512, 1513, 1514, 1515, 1516, 1517+2048
, 1518, 1519, 1520, 1521, 1522, 1523, 1524, 1525, 1526, 1527, 1528+2048
, 1529, 1530, 1531, 1532, 1533, 1534, 1535, 1536, 1537, 1538, 1539+2048
, 1540, 1541, 1542, 1543, 1544, 1545, 1546, 1547, 1548, 1549, 1550+2048
, 1551, 1552, 1553, 1554, 1555, 1556, 1557, 1558, 1559, 1560, 1561+2048
, 1562, 1563, 1564, 1565, 1566, 1567, 1568, 1569, 1570, 1571, 1572+2048
, 1573, 1574, 1575, 1576, 1577, 1578, 1579, 1580, 1581, 1582, 1583+2048

,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9+2048
,   10,   11,   12,   13,   14,   15,   16,   17,   18,   19+2048
,   20,   21,   22,   23,   24,   25,   26,   27,   28,   29+2048
,   30,   31,   32,   33,   34,   35,   36,   37,   38,   39+2048
,   40,   41,   42,   43,   44,   45,   46,   47,   48,   49+2048
,   50,   51,   52,   53,   54,   55,   56,   57,   58,   59+2048
,   60,   61,   62,   63,   64,   65,   66,   67,   68,   69+2048
,   70,   71,   72,   73,   74,   75,   76,   77,   78,   79+2048
,   80,   81,   82,   83,   84,   85,   86,   87,   88,   89+2048
,   90,   91,   92,   93,   94,   95,   96,   97,   98,   99+2048
,  100,  101,  102,  103,  104,  105,  106,  107,  108,  109+2048
,  110,  111,  112,  113,  114,  115,  116,  117,  118,  119+2048
,  120,  121,  122,  123,  124,  125,  126,  127,  128,  129+2048
,  130,  131,  132,  133,  134,  135,  136,  137,  138,  139+2048
,  140,  141,  142,  143,  144,  145,  146,  147,  148,  149+2048
,  150,  151,  152,  153,  154,  155,  156,  157,  158,  159+2048
,  160,  161,  162,  163,  164,  165,  166,  167,  168,  169+2048
,  170,  171,  172,  173,  174,  175,  176,  177,  178,  179+2048
,  180,  181,  182,  183,  184,  185,  186,  187,  188,  189+2048
,  190,  191,  192,  193,  194,  195,  196,  197,  198,  199+2048
,  200,  201,  202,  203,  204,  205,  206,  207,  208,  209+2048
,  210,  211,  212,  213,  214,  215,  216,  217,  218,  219+2048
,  220,  221,  222,  223,  224,  225,  226,  227,  228,  229+2048
,  230,  231,  232,  233,  234,  235,  236,  237,  238,  239+2048
,  240,  241,  242,  243,  244,  245,  246,  247,  248,  249+2048
,  250,  251,  252,  253,  254,  255,  256,  257,  258,  259+2048
,  260,  261,  262,  263,  264,  265,  266,  267,  268,  269+2048
,  270,  271,  272,  273,  274,  275,  276,  277,  278,  279+2048
,  280,  281,  282,  283,  284,  285,  286,  287,  288,  289+2048
,  290,  291,  292,  293,  294,  295,  296,  297,  298,  299+2048
,  300,  301,  302,  303,  304,  305,  306,  307,  308,  309+2048
,  310,  311,  312,  313,  314,  315,  316,  317,  318,  319+2048
,  320,  321,  322,  323,  324,  325,  326,  327,  328,  329+2048
,  330,  331,  332,  333,  334,  335,  336,  337,  338,  339+2048
,  340,  341,  342,  343,  344,  345,  346,  347,  348,  349+2048
,  350,  351,  352,  353,  354,  355,  356,  357,  358,  359+2048
,  360,  361,  362,  363,  364,  365,  366,  367,  368,  369+2048
,  370,  371,  372,  373,  374,  375,  376,  377,  378,  379+2048
,  380,  381,  382,  383,  384,  385,  386,  387,  388,  389+2048
,  390,  391,  392,  393,  394,  395,  396,  397,  398,  399+2048
,  400,  401,  402,  403,  404,  405,  406,  407,  408,  409+2048
,  410,  411,  412,  413,  414,  415,  416,  417,  418,  419+2048
,  420,  421,  422,  423,  424,  425,  426,  427,  428,  429+2048
,  430,  431,  432,  433,  434,  435,  436,  437,  438,  439+2048
,  440,  441,  442,  443,  444,  445,  446,  447,  448,  449+2048
,  450,  451,  452,  453,  454,  455,  456,  457,  458,  459+2048
,  460,  461,  462,  463,  464,  465,  466,  467,  468,  469+2048
,  470,  471,  472,  473,  474,  475,  476,  477,  478,  479+2048
,  480,  481,  482,  483,  484,  485,  486,  487,  488,  489+2048
,  490,  491,  492,  493,  494,  495,  496,  497,  498,  499+2048
,  500,  501,  502,  503,  504,  505,  506,  507,  508,  509+2048
,  510,  511,  512,  513,  514,  515,  516,  517,  518,  519+2048
,  520,  521,  522,  523,  524,  525,  526,  527,  528,  529+2048
,  530,  531,  532,  533,  534,  535,  536,  537,  538,  539+2048
,  540,  541,  542,  543,  544,  545,  546,  547,  548,  549+2048
,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559+2048
,  560,  561,  562,  563,  564,  565,  566,  567,  568,  569+2048
,  570,  571,  572,  573,  574,  575,  576,  577,  578,  579+2048
,  580,  581,  582,  583,  584,  585,  586,  587,  588,  589+2048
,  590,  591,  592,  593,  594,  595,  596,  597,  598,  599+2048
,  600,  601,  602,  603,  604,  605,  606,  607,  608,  609+2048
,  610,  611,  612,  613,  614,  615,  616,  617,  618,  619+2048
,  620,  621,  622,  623,  624,  625,  626,  627,  628,  629+2048
,  630,  631,  632,  633,  634,  635,  636,  637,  638,  639+2048
,  640,  641,  642,  643,  644,  645,  646,  647,  648,  649+2048
,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659+2048
,  660,  661,  662,  663,  664,  665,  666,  667,  668,  669+2048
,  670,  671,  672,  673,  674,  675,  676,  677,  678,  679+2048
,  680,  681,  682,  683,  684,  685,  686,  687,  688,  689+2048
,  690,  691,  692,  693,  694,  695,  696,  697,  698,  699+2048
,  700,  701,  702,  703,  704,  705,  706,  707,  708,  709+2048
,  710,  711,  712,  713,  714,  715,  716,  717,  718,  719+2048
,  720,  721,  722,  723,  724,  725,  726,  727,  728,  729+2048
,  730,  731,  732,  733,  734,  735,  736,  737,  738,  739+2048
,  740,  741,  742,  743,  744,  745,  746,  747,  748,  749+2048
,  750,  751,  752,  753,  754,  755,  756,  757,  758,  759+2048
,  760,  761,  762,  763,  764,  765,  766,  767,  768,  769+2048
,  770,  771,  772,  773,  774,  775,  776,  777,  778,  779+2048
,  780,  781,  782,  783,  784,  785,  786,  787,  788,  789+2048
,  790,  791,  792,  793,  794,  795,  796,  797,  798,  799+2048
,  800,  801,  802,  803,  804,  805,  806,  807,  808,  809+2048
,  810,  811,  812,  813,  814,  815,  816,  817,  818,  819+2048
,  820,  821,  822,  823,  824,  825,  826,  827,  828,  829+2048
,  830,  831,  832,  833,  834,  835,  836,  837,  838,  839+2048
,  840,  841,  842,  843,  844,  845,  846,  847,  848,  849+2048
,  850,  851,  852,  853,  854,  855,  856,  857,  858,  859+2048
,  860,  861,  862,  863,  864,  865,  866,  867,  868,  869+2048
,  870,  871,  872,  873,  874,  875,  876,  877,  878,  879+2048
,  880,  881,  882,  883,  884,  885,  886,  887,  888,  889+2048
,  890,  891,  892,  893,  894,  895,  896,  897,  898,  899+2048
,  900,  901,  902,  903,  904,  905,  906,  907,  908,  909+2048
,  910,  911,  912,  913,  914,  915,  916,  917,  918,  919+2048
,  920,  921,  922,  923,  924,  925,  926,  927,  928,  929+2048
,  930,  931,  932,  933,  934,  935,  936,  937,  938,  939+2048
,  940,  941,  942,  943,  944,  945,  946,  947,  948,  949+2048
,  950,  951,  952,  953,  954,  955,  956,  957,  958,  959+2048
,  960,  961,  962,  963,  964,  965,  966,  967,  968,  969+2048
,  970,  971,  972,  973,  974,  975,  976,  977,  978,  979+2048
,  980,  981,  982,  983,  984,  985,  986,  987,  988,  989+2048
,  990,  991,  992,  993,  994,  995,  996,  997,  998,  999+2048
, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009+2048
, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019+2048
, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029+2048
, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039+2048
, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049+2048
, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059+2048
, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069+2048
, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079+2048
, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089+2048
, 1090, 1091, 1092, 1093, 1094, 1095, 1096, 1097, 1098, 1099+2048
, 1100, 1101, 1102, 1103, 1104, 1105, 1106, 1107, 1108, 1109+2048
, 1110, 1111, 1112, 1113, 1114, 1115, 1116, 1117, 1118, 1119+2048
, 1120, 1121, 1122, 1123, 1124, 1125, 1126, 1127, 1128, 1129+2048
, 1130, 1131, 1132, 1133, 1134, 1135, 1136, 1137, 1138, 1139+2048
, 1140, 1141, 1142, 1143, 1144, 1145, 1146, 1147, 1148, 1149+2048
, 1150, 1151, 1152, 1153, 1154, 1155, 1156, 1157, 1158, 1159+2048
, 1160, 1161, 1162, 1163, 1164, 1165, 1166, 1167, 1168, 1169+2048
, 1170, 1171, 1172, 1173, 1174, 1175, 1176, 1177, 1178, 1179+2048
, 1180, 1181, 1182, 1183, 1184, 1185, 1186, 1187, 1188, 1189+2048
, 1190, 1191, 1192, 1193, 1194, 1195, 1196, 1197, 1198, 1199+2048

,   33,   34,   35,   36,   37,   38,   39,   40,   41+2048
,  165,  166,  167,  168,  169,  170,  171,  172,  173+2048
,  297,  298,  299,  300,  301,  302,  303,  304,  305+2048
,  429,  430,  431,  432,  433,  434,  435,  436,  437+2048
,  561,  562,  563,  564,  565,  566,  567,  568,  569+2048
,  693,  694,  695,  696,  697,  698,  699,  700,  701+2048
,  825,  826,  827,  828,  829,  830,  831,  832,  833+2048
,  957,  958,  959,  960,  961,  962,  963,  964,  965+2048
,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9+2048
,   42,   43,   44,   45,   46,   47,   48,   49,   50,   51+2048
,   99,  100,  101,  102,  103,  104,  105,  106,  107,  108+2048
,  132,  133,  134,  135,  136,  137,  138,  139,  140,  141+2048
,  174,  175,  176,  177,  178,  179,  180,  181,  182,  183+2048
,  231,  232,  233,  234,  235,  236,  237,  238,  239,  240+2048
,  264,  265,  266,  267,  268,  269,  270,  271,  272,  273+2048
,  306,  307,  308,  309,  310,  311,  312,  313,  314,  315+2048
,  363,  364,  365,  366,  367,  368,  369,  370,  371,  372+2048
,  396,  397,  398,  399,  400,  401,  402,  403,  404,  405+2048
,  438,  439,  440,  441,  442,  443,  444,  445,  446,  447+2048
,  495,  496,  497,  498,  499,  500,  501,  502,  503,  504+2048
,  528,  529,  530,  531,  532,  533,  534,  535,  536,  537+2048
,  570,  571,  572,  573,  574,  575,  576,  577,  578,  579+2048
,  627,  628,  629,  630,  631,  632,  633,  634,  635,  636+2048
,  660,  661,  662,  663,  664,  665,  666,  667,  668,  669+2048
,  702,  703,  704,  705,  706,  707,  708,  709,  710,  711+2048
,  759,  760,  761,  762,  763,  764,  765,  766,  767,  768+2048
,  792,  793,  794,  795,  796,  797,  798,  799,  800,  801+2048
,  834,  835,  836,  837,  838,  839,  840,  841,  842,  843+2048
,  891,  892,  893,  894,  895,  896,  897,  898,  899,  900+2048
,  924,  925,  926,  927,  928,  929,  930,  931,  932,  933+2048
,  966,  967,  968,  969,  970,  971,  972,  973,  974,  975+2048
, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032+2048
,   22,   23,   24,   25,   26,   27,   28,   29,   30,   31,   32+2048
,   65,   66,   67,   68,   69,   70,   71,   72,   73,   74,   75+2048
,   88,   89,   90,   91,   92,   93,   94,   95,   96,   97,   98+2048
,  109,  110,  111,  112,  113,  114,  115,  116,  117,  118,  119+2048
,  154,  155,  156,  157,  158,  159,  160,  161,  162,  163,  164+2048
,  197,  198,  199,  200,  201,  202,  203,  204,  205,  206,  207+2048
,  220,  221,  222,  223,  224,  225,  226,  227,  228,  229,  230+2048
,  241,  242,  243,  244,  245,  246,  247,  248,  249,  250,  251+2048
,  286,  287,  288,  289,  290,  291,  292,  293,  294,  295,  296+2048
,  329,  330,  331,  332,  333,  334,  335,  336,  337,  338,  339+2048
,  352,  353,  354,  355,  356,  357,  358,  359,  360,  361,  362+2048
,  373,  374,  375,  376,  377,  378,  379,  380,  381,  382,  383+2048
,  418,  419,  420,  421,  422,  423,  424,  425,  426,  427,  428+2048
,  461,  462,  463,  464,  465,  466,  467,  468,  469,  470,  471+2048
,  484,  485,  486,  487,  488,  489,  490,  491,  492,  493,  494+2048
,  505,  506,  507,  508,  509,  510,  511,  512,  513,  514,  515+2048
,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559,  560+2048
,  593,  594,  595,  596,  597,  598,  599,  600,  601,  602,  603+2048
,  616,  617,  618,  619,  620,  621,  622,  623,  624,  625,  626+2048
,  637,  638,  639,  640,  641,  642,  643,  644,  645,  646,  647+2048
,  682,  683,  684,  685,  686,  687,  688,  689,  690,  691,  692+2048
,  725,  726,  727,  728,  729,  730,  731,  732,  733,  734,  735+2048
,  748,  749,  750,  751,  752,  753,  754,  755,  756,  757,  758+2048
,  769,  770,  771,  772,  773,  774,  775,  776,  777,  778,  779+2048
,  814,  815,  816,  817,  818,  819,  820,  821,  822,  823,  824+2048
,  857,  858,  859,  860,  861,  862,  863,  864,  865,  866,  867+2048
,  880,  881,  882,  883,  884,  885,  886,  887,  888,  889,  890+2048
,  901,  902,  903,  904,  905,  906,  907,  908,  909,  910,  911+2048
,  946,  947,  948,  949,  950,  951,  952,  953,  954,  955,  956+2048
,  989,  990,  991,  992,  993,  994,  995,  996,  997,  998,  999+2048
, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022+2048
, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043+2048
,   10,   11,   12,   13,   14,   15,   16,   17,   18,   19,   20,   21+2048
,   76,   77,   78,   79,   80,   81,   82,   83,   84,   85,   86,   87+2048
,  120,  121,  122,  123,  124,  125,  126,  127,  128,  129,  130,  131+2048
,  142,  143,  144,  145,  146,  147,  148,  149,  150,  151,  152,  153+2048
,  208,  209,  210,  211,  212,  213,  214,  215,  216,  217,  218,  219+2048
,  252,  253,  254,  255,  256,  257,  258,  259,  260,  261,  262,  263+2048
,  274,  275,  276,  277,  278,  279,  280,  281,  282,  283,  284,  285+2048
,  340,  341,  342,  343,  344,  345,  346,  347,  348,  349,  350,  351+2048
,  384,  385,  386,  387,  388,  389,  390,  391,  392,  393,  394,  395+2048
,  406,  407,  408,  409,  410,  411,  412,  413,  414,  415,  416,  417+2048
,  472,  473,  474,  475,  476,  477,  478,  479,  480,  481,  482,  483+2048
,  516,  517,  518,  519,  520,  521,  522,  523,  524,  525,  526,  527+2048
,  538,  539,  540,  541,  542,  543,  544,  545,  546,  547,  548,  549+2048
,  604,  605,  606,  607,  608,  609,  610,  611,  612,  613,  614,  615+2048
,  648,  649,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659+2048
,  670,  671,  672,  673,  674,  675,  676,  677,  678,  679,  680,  681+2048
,  736,  737,  738,  739,  740,  741,  742,  743,  744,  745,  746,  747+2048
,  780,  781,  782,  783,  784,  785,  786,  787,  788,  789,  790,  791+2048
,  802,  803,  804,  805,  806,  807,  808,  809,  810,  811,  812,  813+2048
,  868,  869,  870,  871,  872,  873,  874,  875,  876,  877,  878,  879+2048
,  912,  913,  914,  915,  916,  917,  918,  919,  920,  921,  922,  923+2048
,  934,  935,  936,  937,  938,  939,  940,  941,  942,  943,  944,  945+2048
, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011+2048
, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055+2048
,   52,   53,   54,   55,   56,   57,   58,   59,   60,   61,   62,   63,   64+2048
,  184,  185,  186,  187,  188,  189,  190,  191,  192,  193,  194,  195,  196+2048
,  316,  317,  318,  319,  320,  321,  322,  323,  324,  325,  326,  327,  328+2048
,  448,  449,  450,  451,  452,  453,  454,  455,  456,  457,  458,  459,  460+2048
,  580,  581,  582,  583,  584,  585,  586,  587,  588,  589,  590,  591,  592+2048
,  712,  713,  714,  715,  716,  717,  718,  719,  720,  721,  722,  723,  724+2048
,  844,  845,  846,  847,  848,  849,  850,  851,  852,  853,  854,  855,  856+2048
,  976,  977,  978,  979,  980,  981,  982,  983,  984,  985,  986,  987,  988+2048

,   12,   13,   14,   15,   16,   17,   18,   19,   20,   21,   22+2048
,  137,  138,  139,  140,  141,  142,  143,  144,  145,  146,  147+2048
,  262,  263,  264,  265,  266,  267,  268,  269,  270,  271,  272+2048
,  387,  388,  389,  390,  391,  392,  393,  394,  395,  396,  397+2048
,  512,  513,  514,  515,  516,  517,  518,  519,  520,  521,  522+2048
,  637,  638,  639,  640,  641,  642,  643,  644,  645,  646,  647+2048
,  762,  763,  764,  765,  766,  767,  768,  769,  770,  771,  772+2048
,  887,  888,  889,  890,  891,  892,  893,  894,  895,  896,  897+2048
,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9,   10,   11+2048
,   36,   37,   38,   39,   40,   41,   42,   43,   44,   45,   46,   47+2048
,   48,   49,   50,   51,   52,   53,   54,   55,   56,   57,   58,   59+2048
,  125,  126,  127,  128,  129,  130,  131,  132,  133,  134,  135,  136+2048
,  161,  162,  163,  164,  165,  166,  167,  168,  169,  170,  171,  172+2048
,  173,  174,  175,  176,  177,  178,  179,  180,  181,  182,  183,  184+2048
,  250,  251,  252,  253,  254,  255,  256,  257,  258,  259,  260,  261+2048
,  286,  287,  288,  289,  290,  291,  292,  293,  294,  295,  296,  297+2048
,  298,  299,  300,  301,  302,  303,  304,  305,  306,  307,  308,  309+2048
,  375,  376,  377,  378,  379,  380,  381,  382,  383,  384,  385,  386+2048
,  411,  412,  413,  414,  415,  416,  417,  418,  419,  420,  421,  422+2048
,  423,  424,  425,  426,  427,  428,  429,  430,  431,  432,  433,  434+2048
,  500,  501,  502,  503,  504,  505,  506,  507,  508,  509,  510,  511+2048
,  536,  537,  538,  539,  540,  541,  542,  543,  544,  545,  546,  547+2048
,  548,  549,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559+2048
,  625,  626,  627,  628,  629,  630,  631,  632,  633,  634,  635,  636+2048
,  661,  662,  663,  664,  665,  666,  667,  668,  669,  670,  671,  672+2048
,  673,  674,  675,  676,  677,  678,  679,  680,  681,  682,  683,  684+2048
,  750,  751,  752,  753,  754,  755,  756,  757,  758,  759,  760,  761+2048
,  786,  787,  788,  789,  790,  791,  792,  793,  794,  795,  796,  797+2048
,  798,  799,  800,  801,  802,  803,  804,  805,  806,  807,  808,  809+2048
,  875,  876,  877,  878,  879,  880,  881,  882,  883,  884,  885,  886+2048
,  911,  912,  913,  914,  915,  916,  917,  918,  919,  920,  921,  922+2048
,  923,  924,  925,  926,  927,  928,  929,  930,  931,  932,  933,  934+2048
,   23,   24,   25,   26,   27,   28,   29,   30,   31,   32,   33,   34,   35+2048
,   60,   61,   62,   63,   64,   65,   66,   67,   68,   69,   70,   71,   72+2048
,   73,   74,   75,   76,   77,   78,   79,   80,   81,   82,   83,   84,   85+2048
,   86,   87,   88,   89,   90,   91,   92,   93,   94,   95,   96,   97,   98+2048
,   99,  100,  101,  102,  103,  104,  105,  106,  107,  108,  109,  110,  111+2048
,  112,  113,  114,  115,  116,  117,  118,  119,  120,  121,  122,  123,  124+2048
,  148,  149,  150,  151,  152,  153,  154,  155,  156,  157,  158,  159,  160+2048
,  185,  186,  187,  188,  189,  190,  191,  192,  193,  194,  195,  196,  197+2048
,  198,  199,  200,  201,  202,  203,  204,  205,  206,  207,  208,  209,  210+2048
,  211,  212,  213,  214,  215,  216,  217,  218,  219,  220,  221,  222,  223+2048
,  224,  225,  226,  227,  228,  229,  230,  231,  232,  233,  234,  235,  236+2048
,  237,  238,  239,  240,  241,  242,  243,  244,  245,  246,  247,  248,  249+2048
,  273,  274,  275,  276,  277,  278,  279,  280,  281,  282,  283,  284,  285+2048
,  310,  311,  312,  313,  314,  315,  316,  317,  318,  319,  320,  321,  322+2048
,  323,  324,  325,  326,  327,  328,  329,  330,  331,  332,  333,  334,  335+2048
,  336,  337,  338,  339,  340,  341,  342,  343,  344,  345,  346,  347,  348+2048
,  349,  350,  351,  352,  353,  354,  355,  356,  357,  358,  359,  360,  361+2048
,  362,  363,  364,  365,  366,  367,  368,  369,  370,  371,  372,  373,  374+2048
,  398,  399,  400,  401,  402,  403,  404,  405,  406,  407,  408,  409,  410+2048
,  435,  436,  437,  438,  439,  440,  441,  442,  443,  444,  445,  446,  447+2048
,  448,  449,  450,  451,  452,  453,  454,  455,  456,  457,  458,  459,  460+2048
,  461,  462,  463,  464,  465,  466,  467,  468,  469,  470,  471,  472,  473+2048
,  474,  475,  476,  477,  478,  479,  480,  481,  482,  483,  484,  485,  486+2048
,  487,  488,  489,  490,  491,  492,  493,  494,  495,  496,  497,  498,  499+2048
,  523,  524,  525,  526,  527,  528,  529,  530,  531,  532,  533,  534,  535+2048
,  560,  561,  562,  563,  564,  565,  566,  567,  568,  569,  570,  571,  572+2048
,  573,  574,  575,  576,  577,  578,  579,  580,  581,  582,  583,  584,  585+2048
,  586,  587,  588,  589,  590,  591,  592,  593,  594,  595,  596,  597,  598+2048
,  599,  600,  601,  602,  603,  604,  605,  606,  607,  608,  609,  610,  611+2048
,  612,  613,  614,  615,  616,  617,  618,  619,  620,  621,  622,  623,  624+2048
,  648,  649,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659,  660+2048
,  685,  686,  687,  688,  689,  690,  691,  692,  693,  694,  695,  696,  697+2048
,  698,  699,  700,  701,  702,  703,  704,  705,  706,  707,  708,  709,  710+2048
,  711,  712,  713,  714,  715,  716,  717,  718,  719,  720,  721,  722,  723+2048
,  724,  725,  726,  727,  728,  729,  730,  731,  732,  733,  734,  735,  736+2048
,  737,  738,  739,  740,  741,  742,  743,  744,  745,  746,  747,  748,  749+2048
,  773,  774,  775,  776,  777,  778,  779,  780,  781,  782,  783,  784,  785+2048
,  810,  811,  812,  813,  814,  815,  816,  817,  818,  819,  820,  821,  822+2048
,  823,  824,  825,  826,  827,  828,  829,  830,  831,  832,  833,  834,  835+2048
,  836,  837,  838,  839,  840,  841,  842,  843,  844,  845,  846,  847,  848+2048
,  849,  850,  851,  852,  853,  854,  855,  856,  857,  858,  859,  860,  861+2048
,  862,  863,  864,  865,  866,  867,  868,  869,  870,  871,  872,  873,  874+2048
,  898,  899,  900,  901,  902,  903,  904,  905,  906,  907,  908,  909,  910+2048
,  935,  936,  937,  938,  939,  940,  941,  942,  943,  944,  945,  946,  947+2048
,  948,  949,  950,  951,  952,  953,  954,  955,  956,  957,  958,  959,  960+2048
,  961,  962,  963,  964,  965,  966,  967,  968,  969,  970,  971,  972,  973+2048
,  974,  975,  976,  977,  978,  979,  980,  981,  982,  983,  984,  985,  986+2048
,  987,  988,  989,  990,  991,  992,  993,  994,  995,  996,  997,  998,  999+2048

,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9,   10,   11,   12,   13,   14,   15+2048
,   16,   17,   18,   19,   20,   21,   22,   23,   24,   25,   26,   27,   28,   29,   30,   31+2048
,   32,   33,   34,   35,   36,   37,   38,   39,   40,   41,   42,   43,   44,   45,   46,   47+2048
,   48,   49,   50,   51,   52,   53,   54,   55,   56,   57,   58,   59,   60,   61,   62,   63+2048
,  137,  138,  139,  140,  141,  142,  143,  144,  145,  146,  147,  148,  149,  150,  151,  152+2048
,  153,  154,  155,  156,  157,  158,  159,  160,  161,  162,  163,  164,  165,  166,  167,  168+2048
,  169,  170,  171,  172,  173,  174,  175,  176,  177,  178,  179,  180,  181,  182,  183,  184+2048
,  185,  186,  187,  188,  189,  190,  191,  192,  193,  194,  195,  196,  197,  198,  199,  200+2048
,  274,  275,  276,  277,  278,  279,  280,  281,  282,  283,  284,  285,  286,  287,  288,  289+2048
,  290,  291,  292,  293,  294,  295,  296,  297,  298,  299,  300,  301,  302,  303,  304,  305+2048
,  306,  307,  308,  309,  310,  311,  312,  313,  314,  315,  316,  317,  318,  319,  320,  321+2048
,  322,  323,  324,  325,  326,  327,  328,  329,  330,  331,  332,  333,  334,  335,  336,  337+2048
,  411,  412,  413,  414,  415,  416,  417,  418,  419,  420,  421,  422,  423,  424,  425,  426+2048
,  427,  428,  429,  430,  431,  432,  433,  434,  435,  436,  437,  438,  439,  440,  441,  442+2048
,  443,  444,  445,  446,  447,  448,  449,  450,  451,  452,  453,  454,  455,  456,  457,  458+2048
,  459,  460,  461,  462,  463,  464,  465,  466,  467,  468,  469,  470,  471,  472,  473,  474+2048
,  548,  549,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559,  560,  561,  562,  563+2048
,  564,  565,  566,  567,  568,  569,  570,  571,  572,  573,  574,  575,  576,  577,  578,  579+2048
,  580,  581,  582,  583,  584,  585,  586,  587,  588,  589,  590,  591,  592,  593,  594,  595+2048
,  596,  597,  598,  599,  600,  601,  602,  603,  604,  605,  606,  607,  608,  609,  610,  611+2048
,  685,  686,  687,  688,  689,  690,  691,  692,  693,  694,  695,  696,  697,  698,  699,  700+2048
,  701,  702,  703,  704,  705,  706,  707,  708,  709,  710,  711,  712,  713,  714,  715,  716+2048
,  717,  718,  719,  720,  721,  722,  723,  724,  725,  726,  727,  728,  729,  730,  731,  732+2048
,  733,  734,  735,  736,  737,  738,  739,  740,  741,  742,  743,  744,  745,  746,  747,  748+2048
,  822,  823,  824,  825,  826,  827,  828,  829,  830,  831,  832,  833,  834,  835,  836,  837+2048
,  838,  839,  840,  841,  842,  843,  844,  845,  846,  847,  848,  849,  850,  851,  852,  853+2048
,  854,  855,  856,  857,  858,  859,  860,  861,  862,  863,  864,  865,  866,  867,  868,  869+2048
,  870,  871,  872,  873,  874,  875,  876,  877,  878,  879,  880,  881,  882,  883,  884,  885+2048
,  959,  960,  961,  962,  963,  964,  965,  966,  967,  968,  969,  970,  971,  972,  973,  974+2048
,  975,  976,  977,  978,  979,  980,  981,  982,  983,  984,  985,  986,  987,  988,  989,  990+2048
,  991,  992,  993,  994,  995,  996,  997,  998,  999, 1000, 1001, 1002, 1003, 1004, 1005, 1006+2048
, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022+2048
,  120,  121,  122,  123,  124,  125,  126,  127,  128,  129,  130,  131,  132,  133,  134,  135,  136+2048
,  257,  258,  259,  260,  261,  262,  263,  264,  265,  266,  267,  268,  269,  270,  271,  272,  273+2048
,  394,  395,  396,  397,  398,  399,  400,  401,  402,  403,  404,  405,  406,  407,  408,  409,  410+2048
,  531,  532,  533,  534,  535,  536,  537,  538,  539,  540,  541,  542,  543,  544,  545,  546,  547+2048
,  668,  669,  670,  671,  672,  673,  674,  675,  676,  677,  678,  679,  680,  681,  682,  683,  684+2048
,  805,  806,  807,  808,  809,  810,  811,  812,  813,  814,  815,  816,  817,  818,  819,  820,  821+2048
,  942,  943,  944,  945,  946,  947,  948,  949,  950,  951,  952,  953,  954,  955,  956,  957,  958+2048
, 1079, 1080, 1081, 1082, 1083, 1084, 1085, 1086, 1087, 1088, 1089, 1090, 1091, 1092, 1093, 1094, 1095+2048
,   83,   84,   85,   86,   87,   88,   89,   90,   91,   92,   93,   94,   95,   96,   97,   98,   99,  100+2048
,  220,  221,  222,  223,  224,  225,  226,  227,  228,  229,  230,  231,  232,  233,  234,  235,  236,  237+2048
,  357,  358,  359,  360,  361,  362,  363,  364,  365,  366,  367,  368,  369,  370,  371,  372,  373,  374+2048
,  494,  495,  496,  497,  498,  499,  500,  501,  502,  503,  504,  505,  506,  507,  508,  509,  510,  511+2048
,  631,  632,  633,  634,  635,  636,  637,  638,  639,  640,  641,  642,  643,  644,  645,  646,  647,  648+2048
,  768,  769,  770,  771,  772,  773,  774,  775,  776,  777,  778,  779,  780,  781,  782,  783,  784,  785+2048
,  905,  906,  907,  908,  909,  910,  911,  912,  913,  914,  915,  916,  917,  918,  919,  920,  921,  922+2048
, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052, 1053, 1054, 1055, 1056, 1057, 1058, 1059+2048
,   64,   65,   66,   67,   68,   69,   70,   71,   72,   73,   74,   75,   76,   77,   78,   79,   80,   81,   82+2048
,  101,  102,  103,  104,  105,  106,  107,  108,  109,  110,  111,  112,  113,  114,  115,  116,  117,  118,  119+2048
,  201,  202,  203,  204,  205,  206,  207,  208,  209,  210,  211,  212,  213,  214,  215,  216,  217,  218,  219+2048
,  238,  239,  240,  241,  242,  243,  244,  245,  246,  247,  248,  249,  250,  251,  252,  253,  254,  255,  256+2048
,  338,  339,  340,  341,  342,  343,  344,  345,  346,  347,  348,  349,  350,  351,  352,  353,  354,  355,  356+2048
,  375,  376,  377,  378,  379,  380,  381,  382,  383,  384,  385,  386,  387,  388,  389,  390,  391,  392,  393+2048
,  475,  476,  477,  478,  479,  480,  481,  482,  483,  484,  485,  486,  487,  488,  489,  490,  491,  492,  493+2048
,  512,  513,  514,  515,  516,  517,  518,  519,  520,  521,  522,  523,  524,  525,  526,  527,  528,  529,  530+2048
,  612,  613,  614,  615,  616,  617,  618,  619,  620,  621,  622,  623,  624,  625,  626,  627,  628,  629,  630+2048
,  649,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659,  660,  661,  662,  663,  664,  665,  666,  667+2048
,  749,  750,  751,  752,  753,  754,  755,  756,  757,  758,  759,  760,  761,  762,  763,  764,  765,  766,  767+2048
,  786,  787,  788,  789,  790,  791,  792,  793,  794,  795,  796,  797,  798,  799,  800,  801,  802,  803,  804+2048
,  886,  887,  888,  889,  890,  891,  892,  893,  894,  895,  896,  897,  898,  899,  900,  901,  902,  903,  904+2048
,  923,  924,  925,  926,  927,  928,  929,  930,  931,  932,  933,  934,  935,  936,  937,  938,  939,  940,  941+2048
, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041+2048
, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078+2048

,    0,    1,    2,    3,    4,    5,    6,    7,    8,    9,   10,   11,   12,   13,   14,   15,   16,   17,   18,   19,   20,   21,   22,   23,   24,   25,   26+2048
,   27,   28,   29,   30,   31,   32,   33,   34,   35,   36,   37,   38,   39,   40,   41,   42,   43,   44,   45,   46,   47,   48,   49,   50,   51,   52,   53+2048
,   54,   55,   56,   57,   58,   59,   60,   61,   62,   63,   64,   65,   66,   67,   68,   69,   70,   71,   72,   73,   74,   75,   76,   77,   78,   79,   80+2048
,   81,   82,   83,   84,   85,   86,   87,   88,   89,   90,   91,   92,   93,   94,   95,   96,   97,   98,   99,  100,  101,  102,  103,  104,  105,  106,  107+2048
,  108,  109,  110,  111,  112,  113,  114,  115,  116,  117,  118,  119,  120,  121,  122,  123,  124,  125,  126,  127,  128,  129,  130,  131,  132,  133,  134+2048
,  135,  136,  137,  138,  139,  140,  141,  142,  143,  144,  145,  146,  147,  148,  149,  150,  151,  152,  153,  154,  155,  156,  157,  158,  159,  160,  161+2048
,  162,  163,  164,  165,  166,  167,  168,  169,  170,  171,  172,  173,  174,  175,  176,  177,  178,  179,  180,  181,  182,  183,  184,  185,  186,  187,  188+2048
,  189,  190,  191,  192,  193,  194,  195,  196,  197,  198,  199,  200,  201,  202,  203,  204,  205,  206,  207,  208,  209,  210,  211,  212,  213,  214,  215+2048
,  216,  217,  218,  219,  220,  221,  222,  223,  224,  225,  226,  227,  228,  229,  230,  231,  232,  233,  234,  235,  236,  237,  238,  239,  240,  241,  242+2048
,  243,  244,  245,  246,  247,  248,  249,  250,  251,  252,  253,  254,  255,  256,  257,  258,  259,  260,  261,  262,  263,  264,  265,  266,  267,  268,  269+2048
,  270,  271,  272,  273,  274,  275,  276,  277,  278,  279,  280,  281,  282,  283,  284,  285,  286,  287,  288,  289,  290,  291,  292,  293,  294,  295,  296+2048
,  297,  298,  299,  300,  301,  302,  303,  304,  305,  306,  307,  308,  309,  310,  311,  312,  313,  314,  315,  316,  317,  318,  319,  320,  321,  322,  323+2048
,  324,  325,  326,  327,  328,  329,  330,  331,  332,  333,  334,  335,  336,  337,  338,  339,  340,  341,  342,  343,  344,  345,  346,  347,  348,  349,  350+2048
,  351,  352,  353,  354,  355,  356,  357,  358,  359,  360,  361,  362,  363,  364,  365,  366,  367,  368,  369,  370,  371,  372,  373,  374,  375,  376,  377+2048
,  378,  379,  380,  381,  382,  383,  384,  385,  386,  387,  388,  389,  390,  391,  392,  393,  394,  395,  396,  397,  398,  399,  400,  401,  402,  403,  404+2048
,  405,  406,  407,  408,  409,  410,  411,  412,  413,  414,  415,  416,  417,  418,  419,  420,  421,  422,  423,  424,  425,  426,  427,  428,  429,  430,  431+2048
,  432,  433,  434,  435,  436,  437,  438,  439,  440,  441,  442,  443,  444,  445,  446,  447,  448,  449,  450,  451,  452,  453,  454,  455,  456,  457,  458+2048
,  459,  460,  461,  462,  463,  464,  465,  466,  467,  468,  469,  470,  471,  472,  473,  474,  475,  476,  477,  478,  479,  480,  481,  482,  483,  484,  485+2048
,  486,  487,  488,  489,  490,  491,  492,  493,  494,  495,  496,  497,  498,  499,  500,  501,  502,  503,  504,  505,  506,  507,  508,  509,  510,  511,  512+2048
,  513,  514,  515,  516,  517,  518,  519,  520,  521,  522,  523,  524,  525,  526,  527,  528,  529,  530,  531,  532,  533,  534,  535,  536,  537,  538,  539+2048
,  540,  541,  542,  543,  544,  545,  546,  547,  548,  549,  550,  551,  552,  553,  554,  555,  556,  557,  558,  559,  560,  561,  562,  563,  564,  565,  566+2048
,  567,  568,  569,  570,  571,  572,  573,  574,  575,  576,  577,  578,  579,  580,  581,  582,  583,  584,  585,  586,  587,  588,  589,  590,  591,  592,  593+2048
,  594,  595,  596,  597,  598,  599,  600,  601,  602,  603,  604,  605,  606,  607,  608,  609,  610,  611,  612,  613,  614,  615,  616,  617,  618,  619,  620+2048
,  621,  622,  623,  624,  625,  626,  627,  628,  629,  630,  631,  632,  633,  634,  635,  636,  637,  638,  639,  640,  641,  642,  643,  644,  645,  646,  647+2048
,  648,  649,  650,  651,  652,  653,  654,  655,  656,  657,  658,  659,  660,  661,  662,  663,  664,  665,  666,  667,  668,  669,  670,  671,  672,  673,  674+2048
,  675,  676,  677,  678,  679,  680,  681,  682,  683,  684,  685,  686,  687,  688,  689,  690,  691,  692,  693,  694,  695,  696,  697,  698,  699,  700,  701+2048
,  702,  703,  704,  705,  706,  707,  708,  709,  710,  711,  712,  713,  714,  715,  716,  717,  718,  719,  720,  721,  722,  723,  724,  725,  726,  727,  728+2048
,  729,  730,  731,  732,  733,  734,  735,  736,  737,  738,  739,  740,  741,  742,  743,  744,  745,  746,  747,  748,  749,  750,  751,  752,  753,  754,  755+2048
,  756,  757,  758,  759,  760,  761,  762,  763,  764,  765,  766,  767,  768,  769,  770,  771,  772,  773,  774,  775,  776,  777,  778,  779,  780,  781,  782+2048
,  783,  784,  785,  786,  787,  788,  789,  790,  791,  792,  793,  794,  795,  796,  797,  798,  799,  800,  801,  802,  803,  804,  805,  806,  807,  808,  809+2048
,  810,  811,  812,  813,  814,  815,  816,  817,  818,  819,  820,  821,  822,  823,  824,  825,  826,  827,  828,  829,  830,  831,  832,  833,  834,  835,  836+2048
,  837,  838,  839,  840,  841,  842,  843,  844,  845,  846,  847,  848,  849,  850,  851,  852,  853,  854,  855,  856,  857,  858,  859,  860,  861,  862,  863+2048
,  864,  865,  866,  867,  868,  869,  870,  871,  872,  873,  874,  875,  876,  877,  878,  879,  880,  881,  882,  883,  884,  885,  886,  887,  888,  889,  890+2048
,  891,  892,  893,  894,  895,  896,  897,  898,  899,  900,  901,  902,  903,  904,  905,  906,  907,  908,  909,  910,  911,  912,  913,  914,  915,  916,  917+2048
,  918,  919,  920,  921,  922,  923,  924,  925,  926,  927,  928,  929,  930,  931,  932,  933,  934,  935,  936,  937,  938,  939,  940,  941,  942,  943,  944+2048
,  945,  946,  947,  948,  949,  950,  951,  952,  953,  954,  955,  956,  957,  958,  959,  960,  961,  962,  963,  964,  965,  966,  967,  968,  969,  970,  971+2048
,  972,  973,  974,  975,  976,  977,  978,  979,  980,  981,  982,  983,  984,  985,  986,  987,  988,  989,  990,  991,  992,  993,  994,  995,  996,  997,  998+2048
,  999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019, 1020, 1021, 1022, 1023, 1024, 1025+2048
, 1026, 1027, 1028, 1029, 1030, 1031, 1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043, 1044, 1045, 1046, 1047, 1048, 1049, 1050, 1051, 1052+2048
, 1053, 1054, 1055, 1056, 1057, 1058, 1059, 1060, 1061, 1062, 1063, 1064, 1065, 1066, 1067, 1068, 1069, 1070, 1071, 1072, 1073, 1074, 1075, 1076, 1077, 1078, 1079+2048);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , Do'length );
		end if;
	end process;

end Behavioral;