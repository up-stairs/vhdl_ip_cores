----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:58:54 09/16/2011 
-- Design Name: 
-- Module Name:    EdgeMap - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE STD.TEXTIO.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity EdgeMap is
	port(
		clk						: in  std_logic;
		
		Addr					: in  std_logic_vector(13 downto 0);
		Do						: out std_logic_vector(17 downto 0)
	);
end EdgeMap;

architecture Behavioral of EdgeMap is
	type INT_TYPE is array (0 to 12893) of integer;
	constant EdgeMapMemory : INT_TYPE := (
(2**17)*0+(2**8)*  0+  2, (2**17)*1+(2**8)* 12+ 52, 
(2**17)*0+(2**8)*  5+ 47, (2**17)*1+(2**8)* 12+ 95, 
(2**17)*0+(2**8)*  1+154, (2**17)*1+(2**8)* 10+ 49, 
(2**17)*0+(2**8)* 11+101, (2**17)*1+(2**8)* 16+ 33, 
(2**17)*0+(2**8)*  0+ 23, (2**17)*1+(2**8)*  9+ 69, 
(2**17)*0+(2**8)*  1+112, (2**17)*1+(2**8)*  3+ 83, 
(2**17)*1+(2**8)*  3+121, 
(2**17)*0+(2**8)*  9+156, (2**17)*1+(2**8)* 10+ 54, 
(2**17)*0+(2**8)* 11+107, (2**17)*1+(2**8)* 11+ 60, 
(2**17)*0+(2**8)*  8+ 69, (2**17)*1+(2**8)* 13+150, 
(2**17)*0+(2**8)*  2+ 37, (2**17)*1+(2**8)* 11+150, 
(2**17)*0+(2**8)*  0+ 88, (2**17)*1+(2**8)* 10+ 43, 
(2**17)*0+(2**8)*  3+ 68, (2**17)*1+(2**8)* 17+137, 
(2**17)*1+(2**8)*  2+ 50, 
(2**17)*1+(2**8)*  9+134, 
(2**17)*1+(2**8)*  0+ 67, 
(2**17)*0+(2**8)*  0+  4, (2**17)*1+(2**8)*  1+115, 
(2**17)*0+(2**8)*  1+143, (2**17)*1+(2**8)*  2+155, 
(2**17)*0+(2**8)* 14+151, (2**17)*1+(2**8)* 17+177, 
(2**17)*0+(2**8)* 10+107, (2**17)*1+(2**8)* 13+ 43, 
(2**17)*1+(2**8)*  1+ 69, 
(2**17)*0+(2**8)*  2+ 49, (2**17)*1+(2**8)*  3+145, 
(2**17)*0+(2**8)*  3+ 46, (2**17)*1+(2**8)* 15+167, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*1+(2**8)* 14+ 80, 
(2**17)*0+(2**8)*  2+ 72, (2**17)*1+(2**8)* 10+ 83, 
(2**17)*0+(2**8)*  2+170, (2**17)*1+(2**8)* 12+165, 
(2**17)*1+(2**8)* 10+ 52, 
(2**17)*1+(2**8)*  9+107, 
(2**17)*1+(2**8)* 15+ 19, 
(2**17)*0+(2**8)*  0+174, (2**17)*1+(2**8)* 16+ 59, 
(2**17)*1+(2**8)* 12+148, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*1+(2**8)*  2+ 91, 
(2**17)*0+(2**8)*  3+154, (2**17)*1+(2**8)* 13+109, 
(2**17)*0+(2**8)* 12+129, (2**17)*1+(2**8)* 16+ 86, 
(2**17)*0+(2**8)*  2+121, (2**17)*1+(2**8)*  6+169, 
(2**17)*0+(2**8)*  1+148, (2**17)*1+(2**8)*  3+ 36, 
(2**17)*0+(2**8)*  3+ 51, (2**17)*1+(2**8)*  9+  2, 
(2**17)*0+(2**8)*  3+ 94, (2**17)*1+(2**8)* 14+ 47, 
(2**17)*0+(2**8)*  1+ 48, (2**17)*1+(2**8)* 10+154, 
(2**17)*0+(2**8)*  2+100, (2**17)*1+(2**8)*  7+ 32, 
(2**17)*0+(2**8)*  0+ 68, (2**17)*1+(2**8)*  9+ 23, 
(2**17)*0+(2**8)* 10+112, (2**17)*1+(2**8)* 12+ 83, 
(2**17)*1+(2**8)* 12+121, 
(2**17)*0+(2**8)*  0+155, (2**17)*1+(2**8)*  1+ 53, 
(2**17)*0+(2**8)*  2+106, (2**17)*1+(2**8)*  2+ 59, 
(2**17)*0+(2**8)*  4+149, (2**17)*1+(2**8)* 17+ 69, 
(2**17)*0+(2**8)*  2+149, (2**17)*1+(2**8)* 11+ 37, 
(2**17)*0+(2**8)*  1+ 42, (2**17)*1+(2**8)*  9+ 88, 
(2**17)*0+(2**8)*  8+136, (2**17)*1+(2**8)* 12+ 68, 
(2**17)*1+(2**8)* 11+ 50, 
(2**17)*1+(2**8)*  0+133, 
(2**17)*1+(2**8)*  9+ 67, 
(2**17)*0+(2**8)*  9+  4, (2**17)*1+(2**8)* 10+115, 
(2**17)*0+(2**8)* 10+143, (2**17)*1+(2**8)* 11+155, 
(2**17)*0+(2**8)*  5+150, (2**17)*1+(2**8)*  8+176, 
(2**17)*0+(2**8)*  1+106, (2**17)*1+(2**8)*  4+ 42, 
(2**17)*1+(2**8)* 10+ 69, 
(2**17)*0+(2**8)* 11+ 49, (2**17)*1+(2**8)* 12+145, 
(2**17)*0+(2**8)*  6+166, (2**17)*1+(2**8)* 12+ 46, 
(2**17)*0+(2**8)*  5+ 79, (2**17)*1+(2**8)*  9+ 77, 
(2**17)*0+(2**8)*  1+ 82, (2**17)*1+(2**8)* 11+ 72, 
(2**17)*0+(2**8)*  3+164, (2**17)*1+(2**8)* 11+170, 
(2**17)*1+(2**8)*  1+ 51, 
(2**17)*1+(2**8)*  0+106, 
(2**17)*1+(2**8)*  6+ 18, 
(2**17)*0+(2**8)*  7+ 58, (2**17)*1+(2**8)*  9+174, 
(2**17)*1+(2**8)*  3+147, 
(2**17)*0+(2**8)*  9+ 87, (2**17)*1+(2**8)* 11+ 91, 
(2**17)*0+(2**8)*  4+108, (2**17)*1+(2**8)* 12+154, 
(2**17)*0+(2**8)*  3+128, (2**17)*1+(2**8)*  7+ 85, 
(2**17)*0+(2**8)* 11+121, (2**17)*1+(2**8)* 15+169, 
(2**17)*0+(2**8)* 10+148, (2**17)*1+(2**8)* 12+ 36, 


(2**17)*0+(2**8)*  3+ 64, (2**17)*0+(2**8)* 17+ 72, (2**17)*1+(2**8)* 25+166, 
(2**17)*0+(2**8)* 16+101, (2**17)*0+(2**8)* 19+143, (2**17)*1+(2**8)* 19+ 31, 
(2**17)*0+(2**8)* 15+ 49, (2**17)*0+(2**8)* 19+175, (2**17)*1+(2**8)* 21+120, 
(2**17)*0+(2**8)*  0+112, (2**17)*0+(2**8)*  9+126, (2**17)*1+(2**8)* 18+ 62, 
(2**17)*0+(2**8)* 17+ 19, (2**17)*0+(2**8)* 27+ 29, (2**17)*1+(2**8)* 29+ 56, 
(2**17)*0+(2**8)*  5+ 25, (2**17)*0+(2**8)* 16+ 60, (2**17)*1+(2**8)* 18+104, 
(2**17)*0+(2**8)*  1+ 37, (2**17)*0+(2**8)* 15+ 54, (2**17)*1+(2**8)* 16+107, 
(2**17)*0+(2**8)*  2+169, (2**17)*0+(2**8)* 11+ 45, (2**17)*1+(2**8)* 18+ 47, 
(2**17)*0+(2**8)* 16+150, (2**17)*0+(2**8)* 20+130, (2**17)*1+(2**8)* 28+ 65, 
(2**17)*0+(2**8)* 11+160, (2**17)*0+(2**8)* 17+168, (2**17)*1+(2**8)* 17+ 86, 
(2**17)*0+(2**8)*  8+171, (2**17)*0+(2**8)* 15+ 43, (2**17)*1+(2**8)* 18+ 86, 
(2**17)*0+(2**8)*  1+ 50, (2**17)*0+(2**8)*  2+ 38, (2**17)*1+(2**8)* 22+ 66, 
(2**17)*0+(2**8)*  0+115, (2**17)*0+(2**8)*  1+155, (2**17)*1+(2**8)* 20+ 95, 
(2**17)*0+(2**8)*  0+143, (2**17)*0+(2**8)* 19+ 90, (2**17)*1+(2**8)* 27+115, 
(2**17)*0+(2**8)*  2+  7, (2**17)*0+(2**8)*  8+ 15, (2**17)*1+(2**8)* 26+ 81, 
(2**17)*0+(2**8)*  4+ 25, (2**17)*0+(2**8)* 15+107, (2**17)*1+(2**8)* 17+ 33, 
(2**17)*0+(2**8)*  0+ 69, (2**17)*0+(2**8)*  3+145, (2**17)*1+(2**8)* 19+ 72, 
(2**17)*0+(2**8)*  1+ 49, (2**17)*0+(2**8)* 29+169, (2**17)*1+(2**8)* 29+138, 
(2**17)*0+(2**8)*  1+170, (2**17)*0+(2**8)* 10+ 84, (2**17)*1+(2**8)* 17+167, 
(2**17)*0+(2**8)*  1+ 72, (2**17)*0+(2**8)*  4+ 81, (2**17)*1+(2**8)* 15+ 83, 
(2**17)*0+(2**8)*  3+ 90, (2**17)*0+(2**8)* 19+102, (2**17)*1+(2**8)* 21+114, 
(2**17)*0+(2**8)*  3+ 32, (2**17)*0+(2**8)*  4+ 57, (2**17)*1+(2**8)*  7+121, 
(2**17)*0+(2**8)*  3+ 76, (2**17)*0+(2**8)*  9+ 60, (2**17)*1+(2**8)* 15+ 52, 
(2**17)*0+(2**8)*  2+ 56, (2**17)*0+(2**8)*  3+ 12, (2**17)*1+(2**8)*  6+110, 
(2**17)*0+(2**8)*  2+156, (2**17)*0+(2**8)*  4+123, (2**17)*1+(2**8)* 25+ 76, 
(2**17)*0+(2**8)*  1+ 91, (2**17)*0+(2**8)*  7+ 58, (2**17)*1+(2**8)* 18+127, 
(2**17)*0+(2**8)*  4+ 82, (2**17)*0+(2**8)* 15+  7, (2**17)*1+(2**8)* 17+ 59, 
(2**17)*0+(2**8)* 18+118, (2**17)*0+(2**8)* 27+ 54, (2**17)*1+(2**8)* 28+167, 
(2**17)*0+(2**8)*  1+121, (2**17)*0+(2**8)*  9+156, (2**17)*1+(2**8)* 13+ 79, 
(2**17)*0+(2**8)*  0+148, (2**17)*0+(2**8)*  4+159, (2**17)*1+(2**8)*  8+144, 
(2**17)*0+(2**8)*  2+ 71, (2**17)*0+(2**8)* 10+165, (2**17)*1+(2**8)* 18+ 64, 
(2**17)*0+(2**8)*  1+100, (2**17)*0+(2**8)*  4+142, (2**17)*1+(2**8)*  4+ 30, 
(2**17)*0+(2**8)*  0+ 48, (2**17)*0+(2**8)*  4+174, (2**17)*1+(2**8)*  6+119, 
(2**17)*0+(2**8)*  3+ 61, (2**17)*0+(2**8)* 15+112, (2**17)*1+(2**8)* 24+126, 
(2**17)*0+(2**8)*  2+ 18, (2**17)*0+(2**8)* 12+ 28, (2**17)*1+(2**8)* 14+ 55, 
(2**17)*0+(2**8)*  1+ 59, (2**17)*0+(2**8)*  3+103, (2**17)*1+(2**8)* 20+ 25, 
(2**17)*0+(2**8)*  0+ 53, (2**17)*0+(2**8)*  1+106, (2**17)*1+(2**8)* 16+ 37, 
(2**17)*0+(2**8)*  3+ 46, (2**17)*0+(2**8)* 17+169, (2**17)*1+(2**8)* 26+ 45, 
(2**17)*0+(2**8)*  1+149, (2**17)*0+(2**8)*  5+129, (2**17)*1+(2**8)* 13+ 64, 
(2**17)*0+(2**8)*  2+167, (2**17)*0+(2**8)*  2+ 85, (2**17)*1+(2**8)* 26+160, 
(2**17)*0+(2**8)*  0+ 42, (2**17)*0+(2**8)*  3+ 85, (2**17)*1+(2**8)* 23+171, 
(2**17)*0+(2**8)*  7+ 65, (2**17)*0+(2**8)* 16+ 50, (2**17)*1+(2**8)* 17+ 38, 
(2**17)*0+(2**8)*  5+ 94, (2**17)*0+(2**8)* 15+115, (2**17)*1+(2**8)* 16+155, 
(2**17)*0+(2**8)*  4+ 89, (2**17)*0+(2**8)* 12+114, (2**17)*1+(2**8)* 15+143, 
(2**17)*0+(2**8)* 11+ 80, (2**17)*0+(2**8)* 17+  7, (2**17)*1+(2**8)* 23+ 15, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)*  2+ 32, (2**17)*1+(2**8)* 19+ 25, 
(2**17)*0+(2**8)*  4+ 71, (2**17)*0+(2**8)* 15+ 69, (2**17)*1+(2**8)* 18+145, 
(2**17)*0+(2**8)* 14+168, (2**17)*0+(2**8)* 14+137, (2**17)*1+(2**8)* 16+ 49, 
(2**17)*0+(2**8)*  2+166, (2**17)*0+(2**8)* 16+170, (2**17)*1+(2**8)* 25+ 84, 
(2**17)*0+(2**8)*  0+ 82, (2**17)*0+(2**8)* 16+ 72, (2**17)*1+(2**8)* 19+ 81, 
(2**17)*0+(2**8)*  4+101, (2**17)*0+(2**8)*  6+113, (2**17)*1+(2**8)* 18+ 90, 
(2**17)*0+(2**8)* 18+ 32, (2**17)*0+(2**8)* 19+ 57, (2**17)*1+(2**8)* 22+121, 
(2**17)*0+(2**8)*  0+ 51, (2**17)*0+(2**8)* 18+ 76, (2**17)*1+(2**8)* 24+ 60, 
(2**17)*0+(2**8)* 17+ 56, (2**17)*0+(2**8)* 18+ 12, (2**17)*1+(2**8)* 21+110, 
(2**17)*0+(2**8)* 10+ 75, (2**17)*0+(2**8)* 17+156, (2**17)*1+(2**8)* 19+123, 
(2**17)*0+(2**8)*  3+126, (2**17)*0+(2**8)* 16+ 91, (2**17)*1+(2**8)* 22+ 58, 
(2**17)*0+(2**8)*  0+  6, (2**17)*0+(2**8)*  2+ 58, (2**17)*1+(2**8)* 19+ 82, 
(2**17)*0+(2**8)*  3+117, (2**17)*0+(2**8)* 12+ 53, (2**17)*1+(2**8)* 13+166, 
(2**17)*0+(2**8)* 16+121, (2**17)*0+(2**8)* 24+156, (2**17)*1+(2**8)* 28+ 79, 
(2**17)*0+(2**8)* 15+148, (2**17)*0+(2**8)* 19+159, (2**17)*1+(2**8)* 23+144, 


(2**17)*0+(2**8)*  3+ 82, (2**17)*0+(2**8)*  4+  6, (2**17)*0+(2**8)* 17+165, (2**17)*1+(2**8)* 23+180, 
(2**17)*0+(2**8)*  1+ 93, (2**17)*0+(2**8)*  3+ 70, (2**17)*0+(2**8)*  8+ 86, (2**17)*1+(2**8)* 32+125, 
(2**17)*0+(2**8)*  0+162, (2**17)*0+(2**8)*  5+ 58, (2**17)*0+(2**8)* 13+ 99, (2**17)*1+(2**8)* 23+ 34, 
(2**17)*0+(2**8)*  1+128, (2**17)*0+(2**8)* 20+ 41, (2**17)*0+(2**8)* 20+ 35, (2**17)*1+(2**8)* 32+105, 
(2**17)*0+(2**8)*  3+ 76, (2**17)*0+(2**8)* 24+ 27, (2**17)*0+(2**8)* 26+158, (2**17)*1+(2**8)* 34+ 95, 
(2**17)*0+(2**8)*  4+146, (2**17)*0+(2**8)* 22+109, (2**17)*0+(2**8)* 24+ 31, (2**17)*1+(2**8)* 30+ 92, 
(2**17)*0+(2**8)*  2+166, (2**17)*0+(2**8)*  3+126, (2**17)*0+(2**8)* 13+170, (2**17)*1+(2**8)* 22+119, 
(2**17)*0+(2**8)* 18+105, (2**17)*0+(2**8)* 21+173, (2**17)*0+(2**8)* 23+ 75, (2**17)*1+(2**8)* 30+137, 
(2**17)*0+(2**8)*  9+166, (2**17)*0+(2**8)* 20+114, (2**17)*0+(2**8)* 21+109, (2**17)*1+(2**8)* 22+ 79, 
(2**17)*0+(2**8)*  7+121, (2**17)*0+(2**8)* 10+122, (2**17)*0+(2**8)* 18+ 14, (2**17)*1+(2**8)* 23+ 47, 
(2**17)*0+(2**8)*  0+128, (2**17)*0+(2**8)*  5+ 95, (2**17)*0+(2**8)* 19+  8, (2**17)*1+(2**8)* 35+ 26, 
(2**17)*0+(2**8)*  1+ 31, (2**17)*0+(2**8)*  4+  4, (2**17)*0+(2**8)* 15+ 82, (2**17)*1+(2**8)* 23+ 36, 
(2**17)*0+(2**8)*  9+107, (2**17)*0+(2**8)* 18+ 77, (2**17)*0+(2**8)* 18+ 33, (2**17)*1+(2**8)* 20+164, 
(2**17)*0+(2**8)*  1+ 48, (2**17)*0+(2**8)*  5+ 41, (2**17)*0+(2**8)* 11+ 71, (2**17)*1+(2**8)* 21+ 42, 
(2**17)*0+(2**8)*  5+  9, (2**17)*0+(2**8)* 17+ 49, (2**17)*0+(2**8)* 18+ 12, (2**17)*1+(2**8)* 20+ 36, 
(2**17)*0+(2**8)*  2+ 14, (2**17)*0+(2**8)* 19+ 33, (2**17)*0+(2**8)* 23+173, (2**17)*1+(2**8)* 29+172, 
(2**17)*0+(2**8)*  0+123, (2**17)*0+(2**8)*  2+144, (2**17)*0+(2**8)* 18+ 11, (2**17)*1+(2**8)* 30+161, 
(2**17)*0+(2**8)*  3+140, (2**17)*0+(2**8)*  6+151, (2**17)*0+(2**8)* 10+ 33, (2**17)*1+(2**8)* 21+144, 
(2**17)*0+(2**8)*  3+152, (2**17)*0+(2**8)*  5+ 89, (2**17)*0+(2**8)*  7+ 62, (2**17)*1+(2**8)* 29+ 75, 
(2**17)*0+(2**8)*  4+163, (2**17)*0+(2**8)*  7+ 69, (2**17)*0+(2**8)* 19+104, (2**17)*1+(2**8)* 34+175, 
(2**17)*0+(2**8)*  2+ 33, (2**17)*0+(2**8)* 15+ 83, (2**17)*0+(2**8)* 19+ 16, (2**17)*1+(2**8)* 22+ 81, 
(2**17)*0+(2**8)*  1+ 59, (2**17)*0+(2**8)* 18+ 25, (2**17)*0+(2**8)* 22+179, (2**17)*1+(2**8)* 28+ 82, 
(2**17)*0+(2**8)*  2+134, (2**17)*0+(2**8)*  2+ 16, (2**17)*0+(2**8)*  4+ 88, (2**17)*1+(2**8)* 31+ 37, 
(2**17)*0+(2**8)* 20+ 74, (2**17)*0+(2**8)* 21+100, (2**17)*0+(2**8)* 23+ 15, (2**17)*1+(2**8)* 33+157, 
(2**17)*0+(2**8)*  0+124, (2**17)*0+(2**8)*  1+148, (2**17)*0+(2**8)*  4+ 16, (2**17)*1+(2**8)* 32+167, 
(2**17)*0+(2**8)*  0+149, (2**17)*0+(2**8)*  3+163, (2**17)*0+(2**8)* 26+172, (2**17)*1+(2**8)* 34+136, 
(2**17)*0+(2**8)*  1+105, (2**17)*0+(2**8)* 19+130, (2**17)*0+(2**8)* 22+166, (2**17)*1+(2**8)* 27+137, 
(2**17)*0+(2**8)*  5+179, (2**17)*0+(2**8)* 21+ 82, (2**17)*0+(2**8)* 22+  6, (2**17)*1+(2**8)* 35+165, 
(2**17)*0+(2**8)* 14+124, (2**17)*0+(2**8)* 19+ 93, (2**17)*0+(2**8)* 21+ 70, (2**17)*1+(2**8)* 26+ 86, 
(2**17)*0+(2**8)*  5+ 33, (2**17)*0+(2**8)* 18+162, (2**17)*0+(2**8)* 23+ 58, (2**17)*1+(2**8)* 31+ 99, 
(2**17)*0+(2**8)*  2+ 40, (2**17)*0+(2**8)*  2+ 34, (2**17)*0+(2**8)* 14+104, (2**17)*1+(2**8)* 19+128, 
(2**17)*0+(2**8)*  6+ 26, (2**17)*0+(2**8)*  8+157, (2**17)*0+(2**8)* 16+ 94, (2**17)*1+(2**8)* 21+ 76, 
(2**17)*0+(2**8)*  4+108, (2**17)*0+(2**8)*  6+ 30, (2**17)*0+(2**8)* 12+ 91, (2**17)*1+(2**8)* 22+146, 
(2**17)*0+(2**8)*  4+118, (2**17)*0+(2**8)* 20+166, (2**17)*0+(2**8)* 21+126, (2**17)*1+(2**8)* 31+170, 
(2**17)*0+(2**8)*  0+104, (2**17)*0+(2**8)*  3+172, (2**17)*0+(2**8)*  5+ 74, (2**17)*1+(2**8)* 12+136, 
(2**17)*0+(2**8)*  2+113, (2**17)*0+(2**8)*  3+108, (2**17)*0+(2**8)*  4+ 78, (2**17)*1+(2**8)* 27+166, 
(2**17)*0+(2**8)*  0+ 13, (2**17)*0+(2**8)*  5+ 46, (2**17)*0+(2**8)* 25+121, (2**17)*1+(2**8)* 28+122, 
(2**17)*0+(2**8)*  1+  7, (2**17)*0+(2**8)* 17+ 25, (2**17)*0+(2**8)* 18+128, (2**17)*1+(2**8)* 23+ 95, 
(2**17)*0+(2**8)*  5+ 35, (2**17)*0+(2**8)* 19+ 31, (2**17)*0+(2**8)* 22+  4, (2**17)*1+(2**8)* 33+ 82, 
(2**17)*0+(2**8)*  0+ 76, (2**17)*0+(2**8)*  0+ 32, (2**17)*0+(2**8)*  2+163, (2**17)*1+(2**8)* 27+107, 
(2**17)*0+(2**8)*  3+ 41, (2**17)*0+(2**8)* 19+ 48, (2**17)*0+(2**8)* 23+ 41, (2**17)*1+(2**8)* 29+ 71, 
(2**17)*0+(2**8)*  0+ 11, (2**17)*0+(2**8)*  2+ 35, (2**17)*0+(2**8)* 23+  9, (2**17)*1+(2**8)* 35+ 49, 
(2**17)*0+(2**8)*  1+ 32, (2**17)*0+(2**8)*  5+172, (2**17)*0+(2**8)* 11+171, (2**17)*1+(2**8)* 20+ 14, 
(2**17)*0+(2**8)*  0+ 10, (2**17)*0+(2**8)* 12+160, (2**17)*0+(2**8)* 18+123, (2**17)*1+(2**8)* 20+144, 
(2**17)*0+(2**8)*  3+143, (2**17)*0+(2**8)* 21+140, (2**17)*0+(2**8)* 24+151, (2**17)*1+(2**8)* 28+ 33, 
(2**17)*0+(2**8)* 11+ 74, (2**17)*0+(2**8)* 21+152, (2**17)*0+(2**8)* 23+ 89, (2**17)*1+(2**8)* 25+ 62, 
(2**17)*0+(2**8)*  1+103, (2**17)*0+(2**8)* 16+174, (2**17)*0+(2**8)* 22+163, (2**17)*1+(2**8)* 25+ 69, 
(2**17)*0+(2**8)*  1+ 15, (2**17)*0+(2**8)*  4+ 80, (2**17)*0+(2**8)* 20+ 33, (2**17)*1+(2**8)* 33+ 83, 
(2**17)*0+(2**8)*  0+ 24, (2**17)*0+(2**8)*  4+178, (2**17)*0+(2**8)* 10+ 81, (2**17)*1+(2**8)* 19+ 59, 
(2**17)*0+(2**8)* 13+ 36, (2**17)*0+(2**8)* 20+134, (2**17)*0+(2**8)* 20+ 16, (2**17)*1+(2**8)* 22+ 88, 
(2**17)*0+(2**8)*  2+ 73, (2**17)*0+(2**8)*  3+ 99, (2**17)*0+(2**8)*  5+ 14, (2**17)*1+(2**8)* 15+156, 
(2**17)*0+(2**8)* 14+166, (2**17)*0+(2**8)* 18+124, (2**17)*0+(2**8)* 19+148, (2**17)*1+(2**8)* 22+ 16, 
(2**17)*0+(2**8)*  8+171, (2**17)*0+(2**8)* 16+135, (2**17)*0+(2**8)* 18+149, (2**17)*1+(2**8)* 21+163, 
(2**17)*0+(2**8)*  1+129, (2**17)*0+(2**8)*  4+165, (2**17)*0+(2**8)*  9+136, (2**17)*1+(2**8)* 19+105, 


(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  9+ 77, (2**17)*1+(2**8)* 19+ 69, 
(2**17)*0+(2**8)*  2+114, (2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 21+118, (2**17)*1+(2**8)* 22+ 19, 
(2**17)*0+(2**8)*  3+ 56, (2**17)*0+(2**8)*  4+124, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)* 23+ 72, (2**17)*1+(2**8)* 34+158, 
(2**17)*0+(2**8)*  4+ 40, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 21+127, (2**17)*1+(2**8)* 37+ 61, 
(2**17)*0+(2**8)*  0+127, (2**17)*1+(2**8)*  9+  0, 
(2**17)*0+(2**8)*  6+ 57, (2**17)*0+(2**8)* 10+  0, (2**17)*1+(2**8)* 33+ 62, 
(2**17)*0+(2**8)* 11+  0, (2**17)*1+(2**8)* 13+ 92, 
(2**17)*0+(2**8)*  2+ 70, (2**17)*0+(2**8)* 12+  0, (2**17)*1+(2**8)* 18+ 21, 
(2**17)*0+(2**8)*  0+103, (2**17)*0+(2**8)*  8+ 23, (2**17)*0+(2**8)* 13+  0, (2**17)*1+(2**8)* 34+ 93, 
(2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 25+139, (2**17)*1+(2**8)* 35+ 78, 
(2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 24+ 24, (2**17)*1+(2**8)* 36+179, 
(2**17)*0+(2**8)*  0+ 81, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 19+148, (2**17)*1+(2**8)* 20+ 48, 
(2**17)*0+(2**8)*  0+ 14, (2**17)*0+(2**8)*  0+ 21, (2**17)*0+(2**8)*  7+  4, (2**17)*1+(2**8)* 17+  0, 
(2**17)*0+(2**8)*  4+ 25, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 22+ 49, (2**17)*1+(2**8)* 38+120, 
(2**17)*0+(2**8)* 17+ 15, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 21+ 62, (2**17)*1+(2**8)* 28+ 69, 
(2**17)*0+(2**8)* 22+ 64, (2**17)*0+(2**8)* 24+103, (2**17)*1+(2**8)* 30+  6, 
(2**17)*0+(2**8)*  6+  1, (2**17)*1+(2**8)* 23+ 22, 
(2**17)*0+(2**8)*  3+ 93, (2**17)*0+(2**8)* 11+ 29, (2**17)*0+(2**8)* 24+ 95, (2**17)*1+(2**8)* 32+ 45, 
(2**17)*0+(2**8)* 15+137, (2**17)*0+(2**8)* 21+ 51, (2**17)*1+(2**8)* 22+ 74, 
(2**17)*0+(2**8)*  2+  5, (2**17)*1+(2**8)* 27+134, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  3+ 90, (2**17)*0+(2**8)* 12+156, (2**17)*1+(2**8)* 20+101, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 25+ 81, (2**17)*1+(2**8)* 36+100, 
(2**17)*0+(2**8)*  1+ 96, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  9+ 88, (2**17)*1+(2**8)* 24+130, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)* 21+115, (2**17)*1+(2**8)* 21+ 47, 
(2**17)*0+(2**8)*  3+106, (2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 10+118, (2**17)*0+(2**8)* 23+ 89, (2**17)*1+(2**8)* 31+ 81, 
(2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 29+ 77, (2**17)*1+(2**8)* 39+ 69, 
(2**17)*0+(2**8)*  1+117, (2**17)*0+(2**8)*  2+ 18, (2**17)*0+(2**8)* 22+114, (2**17)*1+(2**8)* 26+  0, 
(2**17)*0+(2**8)*  3+ 71, (2**17)*0+(2**8)* 14+157, (2**17)*0+(2**8)* 23+ 56, (2**17)*0+(2**8)* 24+124, (2**17)*1+(2**8)* 27+  0, 
(2**17)*0+(2**8)*  1+126, (2**17)*0+(2**8)* 17+ 60, (2**17)*0+(2**8)* 24+ 40, (2**17)*1+(2**8)* 28+  0, 
(2**17)*0+(2**8)* 20+127, (2**17)*1+(2**8)* 29+  0, 
(2**17)*0+(2**8)* 13+ 61, (2**17)*0+(2**8)* 26+ 57, (2**17)*1+(2**8)* 30+  0, 
(2**17)*0+(2**8)* 31+  0, (2**17)*1+(2**8)* 33+ 92, 
(2**17)*0+(2**8)* 22+ 70, (2**17)*0+(2**8)* 32+  0, (2**17)*1+(2**8)* 38+ 21, 
(2**17)*0+(2**8)* 14+ 92, (2**17)*0+(2**8)* 20+103, (2**17)*0+(2**8)* 28+ 23, (2**17)*1+(2**8)* 33+  0, 
(2**17)*0+(2**8)*  5+138, (2**17)*0+(2**8)* 15+ 77, (2**17)*1+(2**8)* 34+  0, 
(2**17)*0+(2**8)*  4+ 23, (2**17)*0+(2**8)* 16+178, (2**17)*1+(2**8)* 35+  0, 
(2**17)*0+(2**8)*  0+ 47, (2**17)*0+(2**8)* 20+ 81, (2**17)*0+(2**8)* 36+  0, (2**17)*1+(2**8)* 39+148, 
(2**17)*0+(2**8)* 20+ 14, (2**17)*0+(2**8)* 20+ 21, (2**17)*0+(2**8)* 27+  4, (2**17)*1+(2**8)* 37+  0, 
(2**17)*0+(2**8)*  2+ 48, (2**17)*0+(2**8)* 18+119, (2**17)*0+(2**8)* 24+ 25, (2**17)*1+(2**8)* 38+  0, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*0+(2**8)*  8+ 68, (2**17)*0+(2**8)* 37+ 15, (2**17)*1+(2**8)* 39+  0, 
(2**17)*0+(2**8)*  2+ 63, (2**17)*0+(2**8)*  4+102, (2**17)*1+(2**8)* 10+  5, 
(2**17)*0+(2**8)*  3+ 21, (2**17)*1+(2**8)* 26+  1, 
(2**17)*0+(2**8)*  4+ 94, (2**17)*0+(2**8)* 12+ 44, (2**17)*0+(2**8)* 23+ 93, (2**17)*1+(2**8)* 31+ 29, 
(2**17)*0+(2**8)*  1+ 50, (2**17)*0+(2**8)*  2+ 73, (2**17)*1+(2**8)* 35+137, 
(2**17)*0+(2**8)*  7+133, (2**17)*1+(2**8)* 22+  5, 
(2**17)*0+(2**8)*  0+100, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 23+ 90, (2**17)*1+(2**8)* 32+156, 
(2**17)*0+(2**8)*  5+ 80, (2**17)*0+(2**8)* 16+ 99, (2**17)*1+(2**8)* 21+  0, 
(2**17)*0+(2**8)*  4+129, (2**17)*0+(2**8)* 21+ 96, (2**17)*0+(2**8)* 22+  0, (2**17)*1+(2**8)* 29+ 88, 
(2**17)*0+(2**8)*  1+114, (2**17)*0+(2**8)*  1+ 46, (2**17)*1+(2**8)* 23+  0, 
(2**17)*0+(2**8)*  3+ 88, (2**17)*0+(2**8)* 11+ 80, (2**17)*0+(2**8)* 23+106, (2**17)*0+(2**8)* 24+  0, (2**17)*1+(2**8)* 30+118, 


(2**17)*0+(2**8)*  2+ 86, (2**17)*0+(2**8)*  3+119, (2**17)*0+(2**8)*  6+106, (2**17)*0+(2**8)*  8+ 11, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 27+179, (2**17)*0+(2**8)* 35+ 60, (2**17)*0+(2**8)* 38+ 70, (2**17)*1+(2**8)* 45+136, 
(2**17)*0+(2**8)*  4+ 42, (2**17)*0+(2**8)*  6+161, (2**17)*0+(2**8)*  8+113, (2**17)*0+(2**8)*  9+ 60, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 26+116, (2**17)*0+(2**8)* 28+138, (2**17)*0+(2**8)* 29+180, (2**17)*1+(2**8)* 32+ 56, 
(2**17)*0+(2**8)*  1+ 11, (2**17)*0+(2**8)*  6+ 45, (2**17)*0+(2**8)*  8+157, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 29+176, (2**17)*0+(2**8)* 29+112, (2**17)*0+(2**8)* 35+ 25, (2**17)*0+(2**8)* 43+ 27, (2**17)*1+(2**8)* 52+127, 
(2**17)*0+(2**8)*  1+ 20, (2**17)*0+(2**8)*  2+ 31, (2**17)*0+(2**8)*  4+172, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 22+117, (2**17)*0+(2**8)* 28+156, (2**17)*0+(2**8)* 32+ 86, (2**17)*0+(2**8)* 32+164, (2**17)*1+(2**8)* 37+ 41, 
(2**17)*0+(2**8)*  0+ 15, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 17+158, (2**17)*0+(2**8)* 24+ 94, (2**17)*0+(2**8)* 27+ 61, (2**17)*0+(2**8)* 28+ 35, (2**17)*0+(2**8)* 35+ 79, (2**17)*0+(2**8)* 35+ 50, (2**17)*1+(2**8)* 35+132, 
(2**17)*0+(2**8)*  3+132, (2**17)*0+(2**8)*  7+ 31, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 14+ 48, (2**17)*0+(2**8)* 27+134, (2**17)*0+(2**8)* 28+ 73, (2**17)*0+(2**8)* 30+ 16, (2**17)*0+(2**8)* 31+  2, (2**17)*1+(2**8)* 48+ 81, 
(2**17)*0+(2**8)*  0+ 38, (2**17)*0+(2**8)*  2+147, (2**17)*0+(2**8)*  5+ 74, (2**17)*0+(2**8)*  5+121, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 15+105, (2**17)*0+(2**8)* 34+ 61, (2**17)*0+(2**8)* 35+ 38, (2**17)*1+(2**8)* 50+145, 
(2**17)*0+(2**8)*  2+137, (2**17)*0+(2**8)*  6+ 64, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 19+ 90, (2**17)*0+(2**8)* 27+159, (2**17)*0+(2**8)* 30+ 88, (2**17)*0+(2**8)* 31+117, (2**17)*0+(2**8)* 33+ 23, (2**17)*1+(2**8)* 36+ 74, 
(2**17)*0+(2**8)*  6+153, (2**17)*0+(2**8)* 16+119, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 27+120, (2**17)*0+(2**8)* 32+106, (2**17)*0+(2**8)* 33+ 81, (2**17)*0+(2**8)* 34+157, (2**17)*0+(2**8)* 34+136, (2**17)*1+(2**8)* 48+100, 
(2**17)*0+(2**8)*  4+ 83, (2**17)*0+(2**8)*  5+150, (2**17)*0+(2**8)*  6+ 91, (2**17)*0+(2**8)* 13+166, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 30+116, (2**17)*0+(2**8)* 31+106, (2**17)*0+(2**8)* 32+143, (2**17)*1+(2**8)* 50+131, 
(2**17)*0+(2**8)*  0+ 94, (2**17)*0+(2**8)*  2+173, (2**17)*0+(2**8)*  4+124, (2**17)*0+(2**8)*  7+167, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 22+ 71, (2**17)*0+(2**8)* 30+ 95, (2**17)*0+(2**8)* 32+104, (2**17)*1+(2**8)* 42+ 54, 
(2**17)*0+(2**8)*  3+ 57, (2**17)*0+(2**8)*  6+ 24, (2**17)*0+(2**8)* 12+110, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 20+132, (2**17)*0+(2**8)* 27+ 77, (2**17)*0+(2**8)* 30+ 68, (2**17)*0+(2**8)* 31+ 48, (2**17)*1+(2**8)* 34+ 65, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*0+(2**8)*  1+ 81, (2**17)*0+(2**8)*  3+157, (2**17)*0+(2**8)*  5+177, (2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)* 10+ 38, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 26+136, (2**17)*1+(2**8)* 29+  6, 
(2**17)*0+(2**8)*  1+  7, (2**17)*0+(2**8)*  5+161, (2**17)*0+(2**8)*  7+ 47, (2**17)*0+(2**8)* 12+ 29, (2**17)*0+(2**8)* 20+109, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 28+  6, (2**17)*0+(2**8)* 34+100, (2**17)*1+(2**8)* 35+109, 
(2**17)*0+(2**8)*  2+131, (2**17)*0+(2**8)* 13+168, (2**17)*0+(2**8)* 18+  7, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 27+100, (2**17)*0+(2**8)* 27+ 79, (2**17)*0+(2**8)* 30+110, (2**17)*0+(2**8)* 31+ 12, (2**17)*1+(2**8)* 34+118, 
(2**17)*0+(2**8)*  0+ 21, (2**17)*0+(2**8)*  1+159, (2**17)*0+(2**8)*  6+ 98, (2**17)*0+(2**8)*  7+150, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 30+168, (2**17)*0+(2**8)* 33+ 35, (2**17)*0+(2**8)* 44+ 95, (2**17)*1+(2**8)* 52+142, 
(2**17)*0+(2**8)*  4+ 67, (2**17)*0+(2**8)*  4+ 20, (2**17)*0+(2**8)*  4+131, (2**17)*0+(2**8)* 14+167, (2**17)*0+(2**8)* 24+109, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 29+119, (2**17)*0+(2**8)* 30+176, (2**17)*1+(2**8)* 32+126, 
(2**17)*0+(2**8)*  1+166, (2**17)*0+(2**8)*  2+160, (2**17)*0+(2**8)*  6+ 33, (2**17)*0+(2**8)* 19+136, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 34+  8, (2**17)*0+(2**8)* 35+ 36, (2**17)*0+(2**8)* 35+ 82, (2**17)*1+(2**8)* 38+103, 
(2**17)*0+(2**8)*  0+178, (2**17)*0+(2**8)*  8+ 59, (2**17)*0+(2**8)* 11+ 69, (2**17)*0+(2**8)* 18+135, (2**17)*0+(2**8)* 29+ 86, (2**17)*0+(2**8)* 30+119, (2**17)*0+(2**8)* 33+106, (2**17)*0+(2**8)* 35+ 11, (2**17)*1+(2**8)* 36+  0, 
(2**17)*0+(2**8)*  1+137, (2**17)*0+(2**8)*  2+179, (2**17)*0+(2**8)*  5+ 55, (2**17)*0+(2**8)* 31+ 42, (2**17)*0+(2**8)* 33+161, (2**17)*0+(2**8)* 35+113, (2**17)*0+(2**8)* 36+ 60, (2**17)*0+(2**8)* 37+  0, (2**17)*1+(2**8)* 53+116, 
(2**17)*0+(2**8)*  2+175, (2**17)*0+(2**8)*  2+111, (2**17)*0+(2**8)*  8+ 24, (2**17)*0+(2**8)* 16+ 26, (2**17)*0+(2**8)* 25+126, (2**17)*0+(2**8)* 28+ 11, (2**17)*0+(2**8)* 33+ 45, (2**17)*0+(2**8)* 35+157, (2**17)*1+(2**8)* 38+  0, 
(2**17)*0+(2**8)*  1+155, (2**17)*0+(2**8)*  5+ 85, (2**17)*0+(2**8)*  5+163, (2**17)*0+(2**8)* 10+ 40, (2**17)*0+(2**8)* 28+ 20, (2**17)*0+(2**8)* 29+ 31, (2**17)*0+(2**8)* 31+172, (2**17)*0+(2**8)* 39+  0, (2**17)*1+(2**8)* 49+117, 
(2**17)*0+(2**8)*  0+ 60, (2**17)*0+(2**8)*  1+ 34, (2**17)*0+(2**8)*  8+ 78, (2**17)*0+(2**8)*  8+ 49, (2**17)*0+(2**8)*  8+131, (2**17)*0+(2**8)* 27+ 15, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 44+158, (2**17)*1+(2**8)* 51+ 94, 
(2**17)*0+(2**8)*  0+133, (2**17)*0+(2**8)*  1+ 72, (2**17)*0+(2**8)*  3+ 15, (2**17)*0+(2**8)*  4+  1, (2**17)*0+(2**8)* 21+ 80, (2**17)*0+(2**8)* 30+132, (2**17)*0+(2**8)* 34+ 31, (2**17)*0+(2**8)* 41+  0, (2**17)*1+(2**8)* 41+ 48, 
(2**17)*0+(2**8)*  7+ 60, (2**17)*0+(2**8)*  8+ 37, (2**17)*0+(2**8)* 23+144, (2**17)*0+(2**8)* 27+ 38, (2**17)*0+(2**8)* 29+147, (2**17)*0+(2**8)* 32+ 74, (2**17)*0+(2**8)* 32+121, (2**17)*0+(2**8)* 42+  0, (2**17)*1+(2**8)* 42+105, 
(2**17)*0+(2**8)*  0+158, (2**17)*0+(2**8)*  3+ 87, (2**17)*0+(2**8)*  4+116, (2**17)*0+(2**8)*  6+ 22, (2**17)*0+(2**8)*  9+ 73, (2**17)*0+(2**8)* 29+137, (2**17)*0+(2**8)* 33+ 64, (2**17)*0+(2**8)* 43+  0, (2**17)*1+(2**8)* 46+ 90, 
(2**17)*0+(2**8)*  0+119, (2**17)*0+(2**8)*  5+105, (2**17)*0+(2**8)*  6+ 80, (2**17)*0+(2**8)*  7+156, (2**17)*0+(2**8)*  7+135, (2**17)*0+(2**8)* 21+ 99, (2**17)*0+(2**8)* 33+153, (2**17)*0+(2**8)* 43+119, (2**17)*1+(2**8)* 44+  0, 
(2**17)*0+(2**8)*  3+115, (2**17)*0+(2**8)*  4+105, (2**17)*0+(2**8)*  5+142, (2**17)*0+(2**8)* 23+130, (2**17)*0+(2**8)* 31+ 83, (2**17)*0+(2**8)* 32+150, (2**17)*0+(2**8)* 33+ 91, (2**17)*0+(2**8)* 40+166, (2**17)*1+(2**8)* 45+  0, 
(2**17)*0+(2**8)*  3+ 94, (2**17)*0+(2**8)*  5+103, (2**17)*0+(2**8)* 15+ 53, (2**17)*0+(2**8)* 27+ 94, (2**17)*0+(2**8)* 29+173, (2**17)*0+(2**8)* 31+124, (2**17)*0+(2**8)* 34+167, (2**17)*0+(2**8)* 46+  0, (2**17)*1+(2**8)* 49+ 71, 
(2**17)*0+(2**8)*  0+ 76, (2**17)*0+(2**8)*  3+ 67, (2**17)*0+(2**8)*  4+ 47, (2**17)*0+(2**8)*  7+ 64, (2**17)*0+(2**8)* 30+ 57, (2**17)*0+(2**8)* 33+ 24, (2**17)*0+(2**8)* 39+110, (2**17)*0+(2**8)* 47+  0, (2**17)*1+(2**8)* 47+132, 
(2**17)*0+(2**8)*  2+  5, (2**17)*0+(2**8)* 28+ 61, (2**17)*0+(2**8)* 28+ 81, (2**17)*0+(2**8)* 30+157, (2**17)*0+(2**8)* 32+177, (2**17)*0+(2**8)* 34+ 51, (2**17)*0+(2**8)* 37+ 38, (2**17)*0+(2**8)* 48+  0, (2**17)*1+(2**8)* 53+136, 
(2**17)*0+(2**8)*  1+  5, (2**17)*0+(2**8)*  7+ 99, (2**17)*0+(2**8)*  8+108, (2**17)*0+(2**8)* 28+  7, (2**17)*0+(2**8)* 32+161, (2**17)*0+(2**8)* 34+ 47, (2**17)*0+(2**8)* 39+ 29, (2**17)*0+(2**8)* 47+109, (2**17)*1+(2**8)* 49+  0, 
(2**17)*0+(2**8)*  0+ 99, (2**17)*0+(2**8)*  0+ 78, (2**17)*0+(2**8)*  3+109, (2**17)*0+(2**8)*  4+ 11, (2**17)*0+(2**8)*  7+117, (2**17)*0+(2**8)* 29+131, (2**17)*0+(2**8)* 40+168, (2**17)*0+(2**8)* 45+  7, (2**17)*1+(2**8)* 50+  0, 
(2**17)*0+(2**8)*  3+167, (2**17)*0+(2**8)*  6+ 34, (2**17)*0+(2**8)* 17+ 94, (2**17)*0+(2**8)* 25+141, (2**17)*0+(2**8)* 27+ 21, (2**17)*0+(2**8)* 28+159, (2**17)*0+(2**8)* 33+ 98, (2**17)*0+(2**8)* 34+150, (2**17)*1+(2**8)* 51+  0, 
(2**17)*0+(2**8)*  2+118, (2**17)*0+(2**8)*  3+175, (2**17)*0+(2**8)*  5+125, (2**17)*0+(2**8)* 31+ 67, (2**17)*0+(2**8)* 31+ 20, (2**17)*0+(2**8)* 31+131, (2**17)*0+(2**8)* 41+167, (2**17)*0+(2**8)* 51+109, (2**17)*1+(2**8)* 52+  0, 
(2**17)*0+(2**8)*  7+  7, (2**17)*0+(2**8)*  8+ 35, (2**17)*0+(2**8)*  8+ 81, (2**17)*0+(2**8)* 11+102, (2**17)*0+(2**8)* 28+166, (2**17)*0+(2**8)* 29+160, (2**17)*0+(2**8)* 33+ 33, (2**17)*0+(2**8)* 46+136, (2**17)*1+(2**8)* 53+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  0+154, (2**17)*0+(2**8)*  1+ 96, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 23+ 52, (2**17)*0+(2**8)* 41+ 95, (2**17)*0+(2**8)* 41+ 24, (2**17)*1+(2**8)* 48+ 34, 
(2**17)*0+(2**8)*  0+115, (2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 30+107, (2**17)*0+(2**8)* 31+ 51, (2**17)*0+(2**8)* 40+154, (2**17)*0+(2**8)* 45+ 85, (2**17)*1+(2**8)* 52+  8, 
(2**17)*0+(2**8)*  1+  4, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 31+ 62, (2**17)*0+(2**8)* 32+  4, (2**17)*0+(2**8)* 34+ 72, (2**17)*0+(2**8)* 49+171, (2**17)*1+(2**8)* 51+ 12, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  7+  8, (2**17)*0+(2**8)* 14+ 58, (2**17)*0+(2**8)* 16+ 86, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 30+ 52, (2**17)*0+(2**8)* 31+104, (2**17)*1+(2**8)* 55+ 98, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 28+ 56, (2**17)*0+(2**8)* 31+127, (2**17)*0+(2**8)* 31+118, (2**17)*0+(2**8)* 32+  9, (2**17)*0+(2**8)* 33+118, (2**17)*1+(2**8)* 59+ 38, 
(2**17)*0+(2**8)*  2+104, (2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 27+ 21, (2**17)*0+(2**8)* 30+ 49, (2**17)*0+(2**8)* 35+ 63, (2**17)*0+(2**8)* 36+164, (2**17)*1+(2**8)* 54+ 55, 
(2**17)*0+(2**8)*  2+133, (2**17)*0+(2**8)*  5+161, (2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 12+114, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 22+143, (2**17)*0+(2**8)* 30+ 83, (2**17)*1+(2**8)* 58+  8, 
(2**17)*0+(2**8)*  0+143, (2**17)*0+(2**8)*  2+176, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  9+ 72, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 23+ 16, (2**17)*0+(2**8)* 39+ 84, (2**17)*1+(2**8)* 49+174, 
(2**17)*0+(2**8)*  1+145, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 13+128, (2**17)*0+(2**8)* 18+147, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 30+ 54, (2**17)*0+(2**8)* 32+128, (2**17)*1+(2**8)* 56+ 19, 
(2**17)*0+(2**8)*  0+112, (2**17)*0+(2**8)*  2+113, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 32+ 29, (2**17)*0+(2**8)* 36+129, (2**17)*0+(2**8)* 56+ 79, (2**17)*1+(2**8)* 59+130, 
(2**17)*0+(2**8)*  2+ 88, (2**17)*0+(2**8)*  2+ 78, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 14+ 45, (2**17)*0+(2**8)* 16+ 39, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 42+ 79, (2**17)*1+(2**8)* 50+ 72, 
(2**17)*0+(2**8)*  1+ 32, (2**17)*0+(2**8)*  8+100, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 30+ 43, (2**17)*0+(2**8)* 38+ 48, (2**17)*0+(2**8)* 51+ 90, (2**17)*1+(2**8)* 54+131, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*0+(2**8)*  3+ 11, (2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 17+ 51, (2**17)*0+(2**8)* 20+ 97, (2**17)*0+(2**8)* 27+  0, (2**17)*1+(2**8)* 31+ 47, 
(2**17)*0+(2**8)*  1+ 12, (2**17)*0+(2**8)* 10+ 33, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 15+  5, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 31+115, (2**17)*0+(2**8)* 34+140, (2**17)*1+(2**8)* 57+ 23, 
(2**17)*0+(2**8)*  0+ 69, (2**17)*0+(2**8)*  2+  5, (2**17)*0+(2**8)* 13+ 82, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 32+ 31, (2**17)*0+(2**8)* 47+ 17, (2**17)*1+(2**8)* 55+  5, 
(2**17)*0+(2**8)* 11+ 94, (2**17)*0+(2**8)* 11+ 23, (2**17)*0+(2**8)* 18+ 33, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 30+154, (2**17)*0+(2**8)* 31+ 96, (2**17)*0+(2**8)* 45+  0, (2**17)*1+(2**8)* 53+ 52, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)*  1+ 50, (2**17)*0+(2**8)* 10+153, (2**17)*0+(2**8)* 15+ 84, (2**17)*0+(2**8)* 22+  7, (2**17)*0+(2**8)* 30+115, (2**17)*0+(2**8)* 31+  0, (2**17)*1+(2**8)* 46+  0, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*0+(2**8)*  2+  3, (2**17)*0+(2**8)*  4+ 71, (2**17)*0+(2**8)* 19+170, (2**17)*0+(2**8)* 21+ 11, (2**17)*0+(2**8)* 31+  4, (2**17)*0+(2**8)* 32+  0, (2**17)*1+(2**8)* 47+  0, 
(2**17)*0+(2**8)*  0+ 51, (2**17)*0+(2**8)*  1+103, (2**17)*0+(2**8)* 25+ 97, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 37+  8, (2**17)*0+(2**8)* 44+ 58, (2**17)*0+(2**8)* 46+ 86, (2**17)*1+(2**8)* 48+  0, 
(2**17)*0+(2**8)*  1+126, (2**17)*0+(2**8)*  1+117, (2**17)*0+(2**8)*  2+  8, (2**17)*0+(2**8)*  3+117, (2**17)*0+(2**8)* 29+ 37, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 49+  0, (2**17)*1+(2**8)* 58+ 56, 
(2**17)*0+(2**8)*  0+ 48, (2**17)*0+(2**8)*  5+ 62, (2**17)*0+(2**8)*  6+163, (2**17)*0+(2**8)* 24+ 54, (2**17)*0+(2**8)* 32+104, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 50+  0, (2**17)*1+(2**8)* 57+ 21, 
(2**17)*0+(2**8)*  0+ 82, (2**17)*0+(2**8)* 28+  7, (2**17)*0+(2**8)* 32+133, (2**17)*0+(2**8)* 35+161, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 42+114, (2**17)*0+(2**8)* 51+  0, (2**17)*1+(2**8)* 52+143, 
(2**17)*0+(2**8)*  9+ 83, (2**17)*0+(2**8)* 19+173, (2**17)*0+(2**8)* 30+143, (2**17)*0+(2**8)* 32+176, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 39+ 72, (2**17)*0+(2**8)* 52+  0, (2**17)*1+(2**8)* 53+ 16, 
(2**17)*0+(2**8)*  0+ 53, (2**17)*0+(2**8)*  2+127, (2**17)*0+(2**8)* 26+ 18, (2**17)*0+(2**8)* 31+145, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 43+128, (2**17)*0+(2**8)* 48+147, (2**17)*1+(2**8)* 53+  0, 
(2**17)*0+(2**8)*  2+ 28, (2**17)*0+(2**8)*  6+128, (2**17)*0+(2**8)* 26+ 78, (2**17)*0+(2**8)* 29+129, (2**17)*0+(2**8)* 30+112, (2**17)*0+(2**8)* 32+113, (2**17)*0+(2**8)* 39+  0, (2**17)*1+(2**8)* 54+  0, 
(2**17)*0+(2**8)* 12+ 78, (2**17)*0+(2**8)* 20+ 71, (2**17)*0+(2**8)* 32+ 88, (2**17)*0+(2**8)* 32+ 78, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 44+ 45, (2**17)*0+(2**8)* 46+ 39, (2**17)*1+(2**8)* 55+  0, 
(2**17)*0+(2**8)*  0+ 42, (2**17)*0+(2**8)*  8+ 47, (2**17)*0+(2**8)* 21+ 89, (2**17)*0+(2**8)* 24+130, (2**17)*0+(2**8)* 31+ 32, (2**17)*0+(2**8)* 38+100, (2**17)*0+(2**8)* 41+  0, (2**17)*1+(2**8)* 56+  0, 
(2**17)*0+(2**8)*  1+ 46, (2**17)*0+(2**8)* 30+ 87, (2**17)*0+(2**8)* 33+ 11, (2**17)*0+(2**8)* 37+ 51, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 47+ 51, (2**17)*0+(2**8)* 50+ 97, (2**17)*1+(2**8)* 57+  0, 
(2**17)*0+(2**8)*  1+114, (2**17)*0+(2**8)*  4+139, (2**17)*0+(2**8)* 27+ 22, (2**17)*0+(2**8)* 31+ 12, (2**17)*0+(2**8)* 40+ 33, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 45+  5, (2**17)*1+(2**8)* 58+  0, 
(2**17)*0+(2**8)*  2+ 30, (2**17)*0+(2**8)* 17+ 16, (2**17)*0+(2**8)* 25+  4, (2**17)*0+(2**8)* 30+ 69, (2**17)*0+(2**8)* 32+  5, (2**17)*0+(2**8)* 43+ 82, (2**17)*0+(2**8)* 44+  0, (2**17)*1+(2**8)* 59+  0, 


(2**17)*0+(2**8)*  0+109, (2**17)*0+(2**8)*  8+ 41, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 32+117, (2**17)*0+(2**8)* 44+ 72, (2**17)*0+(2**8)* 45+  6, (2**17)*1+(2**8)* 60+106, 
(2**17)*0+(2**8)*  0+ 42, (2**17)*0+(2**8)*  0+ 75, (2**17)*0+(2**8)*  5+172, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 17+ 81, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 25+140, (2**17)*0+(2**8)* 36+141, (2**17)*0+(2**8)* 53+173, (2**17)*1+(2**8)* 57+ 42, 
(2**17)*0+(2**8)*  0+ 23, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 26+ 41, (2**17)*0+(2**8)* 29+ 54, (2**17)*0+(2**8)* 37+160, (2**17)*0+(2**8)* 40+ 45, (2**17)*0+(2**8)* 46+ 27, (2**17)*1+(2**8)* 49+ 23, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)* 10+125, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 47+144, (2**17)*0+(2**8)* 57+163, (2**17)*1+(2**8)* 63+ 26, 
(2**17)*0+(2**8)*  0+ 80, (2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 18+ 81, (2**17)*0+(2**8)* 18+ 17, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 64+ 69, (2**17)*1+(2**8)* 64+130, 
(2**17)*0+(2**8)*  0+143, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 12+155, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 28+100, (2**17)*0+(2**8)* 33+ 62, (2**17)*0+(2**8)* 34+112, (2**17)*0+(2**8)* 37+144, (2**17)*0+(2**8)* 46+ 76, (2**17)*1+(2**8)* 56+ 30, 
(2**17)*0+(2**8)*  0+133, (2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  6+114, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 19+ 93, (2**17)*0+(2**8)* 26+ 46, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 30+  7, (2**17)*1+(2**8)* 42+ 61, 
(2**17)*0+(2**8)*  0+175, (2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)*  8+ 93, (2**17)*0+(2**8)*  9+126, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 17+ 42, (2**17)*0+(2**8)* 21+128, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 35+168, (2**17)*1+(2**8)* 58+ 97, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  6+174, (2**17)*0+(2**8)* 10+ 55, (2**17)*0+(2**8)* 15+151, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 21+103, (2**17)*0+(2**8)* 22+ 45, (2**17)*0+(2**8)* 29+  0, (2**17)*1+(2**8)* 38+ 86, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 11+ 47, (2**17)*0+(2**8)* 15+ 52, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 29+ 78, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 36+110, (2**17)*1+(2**8)* 55+126, 
(2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  7+164, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 28+ 70, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 33+ 20, (2**17)*0+(2**8)* 47+ 74, (2**17)*0+(2**8)* 49+154, (2**17)*1+(2**8)* 60+  6, 
(2**17)*0+(2**8)*  0+ 28, (2**17)*0+(2**8)*  2+129, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 19+ 41, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 20+ 79, (2**17)*0+(2**8)* 23+ 57, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 34+ 89, (2**17)*1+(2**8)* 65+ 59, 
(2**17)*0+(2**8)* 11+ 71, (2**17)*0+(2**8)* 12+  5, (2**17)*0+(2**8)* 27+105, (2**17)*0+(2**8)* 33+109, (2**17)*0+(2**8)* 41+ 41, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 54+  0, (2**17)*1+(2**8)* 65+117, 
(2**17)*0+(2**8)*  3+140, (2**17)*0+(2**8)* 20+172, (2**17)*0+(2**8)* 24+ 41, (2**17)*0+(2**8)* 33+ 42, (2**17)*0+(2**8)* 33+ 75, (2**17)*0+(2**8)* 38+172, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 50+ 81, (2**17)*0+(2**8)* 55+  0, (2**17)*1+(2**8)* 58+140, 
(2**17)*0+(2**8)*  4+159, (2**17)*0+(2**8)*  7+ 44, (2**17)*0+(2**8)* 13+ 26, (2**17)*0+(2**8)* 16+ 22, (2**17)*0+(2**8)* 33+ 23, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 59+ 41, (2**17)*1+(2**8)* 62+ 54, 
(2**17)*0+(2**8)* 14+143, (2**17)*0+(2**8)* 24+162, (2**17)*0+(2**8)* 30+ 25, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 43+125, (2**17)*0+(2**8)* 45+  0, (2**17)*1+(2**8)* 57+  0, 
(2**17)*0+(2**8)* 31+ 68, (2**17)*0+(2**8)* 31+129, (2**17)*0+(2**8)* 33+ 80, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 51+ 81, (2**17)*0+(2**8)* 51+ 17, (2**17)*1+(2**8)* 58+  0, 
(2**17)*0+(2**8)*  0+ 61, (2**17)*0+(2**8)*  1+111, (2**17)*0+(2**8)*  4+143, (2**17)*0+(2**8)* 13+ 75, (2**17)*0+(2**8)* 23+ 29, (2**17)*0+(2**8)* 33+143, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 45+155, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 59+  0, (2**17)*1+(2**8)* 61+100, 
(2**17)*0+(2**8)*  9+ 60, (2**17)*0+(2**8)* 33+133, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 39+114, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 52+ 93, (2**17)*0+(2**8)* 59+ 46, (2**17)*0+(2**8)* 60+  0, (2**17)*1+(2**8)* 63+  7, 
(2**17)*0+(2**8)*  2+167, (2**17)*0+(2**8)* 25+ 96, (2**17)*0+(2**8)* 33+175, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 41+ 93, (2**17)*0+(2**8)* 42+126, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 50+ 42, (2**17)*0+(2**8)* 54+128, (2**17)*1+(2**8)* 61+  0, 
(2**17)*0+(2**8)*  5+ 85, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 39+174, (2**17)*0+(2**8)* 43+ 55, (2**17)*0+(2**8)* 48+151, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 54+103, (2**17)*0+(2**8)* 55+ 45, (2**17)*1+(2**8)* 62+  0, 
(2**17)*0+(2**8)*  3+109, (2**17)*0+(2**8)* 22+125, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 44+ 47, (2**17)*0+(2**8)* 48+ 52, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 62+ 78, (2**17)*1+(2**8)* 63+  0, 
(2**17)*0+(2**8)*  0+ 19, (2**17)*0+(2**8)* 14+ 73, (2**17)*0+(2**8)* 16+153, (2**17)*0+(2**8)* 27+  5, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 40+164, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 61+ 70, (2**17)*1+(2**8)* 64+  0, 
(2**17)*0+(2**8)*  1+ 88, (2**17)*0+(2**8)* 32+ 58, (2**17)*0+(2**8)* 33+ 28, (2**17)*0+(2**8)* 35+129, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 52+ 41, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 53+ 79, (2**17)*0+(2**8)* 56+ 57, (2**17)*1+(2**8)* 65+  0, 


(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 16+ 90, (2**17)*0+(2**8)* 16+164, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 31+173, (2**17)*0+(2**8)* 37+161, (2**17)*0+(2**8)* 41+ 12, (2**17)*0+(2**8)* 45+106, (2**17)*1+(2**8)* 62+ 81, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 14+ 71, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 22+  6, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 26+ 94, (2**17)*0+(2**8)* 27+135, (2**17)*0+(2**8)* 47+ 48, (2**17)*1+(2**8)* 52+ 17, 
(2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  9+ 43, (2**17)*0+(2**8)* 13+177, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 25+ 36, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 37+ 11, (2**17)*0+(2**8)* 39+ 31, (2**17)*0+(2**8)* 50+114, (2**17)*0+(2**8)* 53+128, (2**17)*1+(2**8)* 63+ 87, 
(2**17)*0+(2**8)*  5+133, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)*  8+ 14, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 20+ 69, (2**17)*0+(2**8)* 20+ 17, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 28+164, (2**17)*0+(2**8)* 30+ 12, (2**17)*1+(2**8)* 36+125, 
(2**17)*0+(2**8)*  1+  9, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 25+ 79, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 42+140, (2**17)*0+(2**8)* 46+102, (2**17)*0+(2**8)* 56+  5, (2**17)*0+(2**8)* 58+139, (2**17)*1+(2**8)* 65+154, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  0+ 78, (2**17)*0+(2**8)*  7+101, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 18+ 23, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 31+ 47, (2**17)*0+(2**8)* 34+177, (2**17)*0+(2**8)* 41+135, (2**17)*1+(2**8)* 59+ 93, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 11+114, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 32+ 87, (2**17)*0+(2**8)* 33+ 28, (2**17)*0+(2**8)* 35+ 45, (2**17)*0+(2**8)* 45+ 19, (2**17)*0+(2**8)* 56+ 12, (2**17)*1+(2**8)* 59+106, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  3+ 36, (2**17)*0+(2**8)*  5+ 97, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 14+ 15, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 26+138, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 33+ 71, (2**17)*0+(2**8)* 50+ 60, (2**17)*1+(2**8)* 58+ 75, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  4+171, (2**17)*0+(2**8)* 12+103, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 13+155, (2**17)*0+(2**8)* 17+115, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 29+  8, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 34+ 58, (2**17)*1+(2**8)* 54+ 52, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)*  9+144, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 32+102, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 38+ 67, (2**17)*0+(2**8)* 43+152, (2**17)*0+(2**8)* 54+124, (2**17)*0+(2**8)* 57+131, (2**17)*1+(2**8)* 64+ 55, 
(2**17)*0+(2**8)*  2+160, (2**17)*0+(2**8)*  6+ 11, (2**17)*0+(2**8)* 10+105, (2**17)*0+(2**8)* 27+ 80, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 51+ 90, (2**17)*0+(2**8)* 51+164, (2**17)*0+(2**8)* 60+  0, (2**17)*1+(2**8)* 66+173, 
(2**17)*0+(2**8)* 12+ 47, (2**17)*0+(2**8)* 17+ 16, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 49+ 71, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 57+  6, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 61+ 94, (2**17)*1+(2**8)* 62+135, 
(2**17)*0+(2**8)*  2+ 10, (2**17)*0+(2**8)*  4+ 30, (2**17)*0+(2**8)* 15+113, (2**17)*0+(2**8)* 18+127, (2**17)*0+(2**8)* 28+ 86, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 44+ 43, (2**17)*0+(2**8)* 48+177, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 60+ 36, (2**17)*1+(2**8)* 62+  0, 
(2**17)*0+(2**8)*  1+124, (2**17)*0+(2**8)* 40+133, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 43+ 14, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 55+ 69, (2**17)*0+(2**8)* 55+ 17, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 63+164, (2**17)*1+(2**8)* 65+ 12, 
(2**17)*0+(2**8)*  7+139, (2**17)*0+(2**8)* 11+101, (2**17)*0+(2**8)* 21+  4, (2**17)*0+(2**8)* 23+138, (2**17)*0+(2**8)* 30+153, (2**17)*0+(2**8)* 36+  9, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 60+ 79, (2**17)*1+(2**8)* 64+  0, 
(2**17)*0+(2**8)*  6+134, (2**17)*0+(2**8)* 24+ 92, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 35+ 78, (2**17)*0+(2**8)* 42+101, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 53+ 23, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 66+ 47, (2**17)*1+(2**8)* 69+177, 
(2**17)*0+(2**8)*  0+ 44, (2**17)*0+(2**8)* 10+ 18, (2**17)*0+(2**8)* 21+ 11, (2**17)*0+(2**8)* 24+105, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 46+114, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 67+ 87, (2**17)*1+(2**8)* 68+ 28, 
(2**17)*0+(2**8)* 15+ 59, (2**17)*0+(2**8)* 23+ 74, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 38+ 36, (2**17)*0+(2**8)* 40+ 97, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 49+ 15, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 61+138, (2**17)*0+(2**8)* 67+  0, (2**17)*1+(2**8)* 68+ 71, 
(2**17)*0+(2**8)* 19+ 51, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 39+171, (2**17)*0+(2**8)* 47+103, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 48+155, (2**17)*0+(2**8)* 52+115, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 64+  8, (2**17)*0+(2**8)* 68+  0, (2**17)*1+(2**8)* 69+ 58, 
(2**17)*0+(2**8)*  3+ 66, (2**17)*0+(2**8)*  8+151, (2**17)*0+(2**8)* 19+123, (2**17)*0+(2**8)* 22+130, (2**17)*0+(2**8)* 29+ 54, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 44+144, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 67+102, (2**17)*1+(2**8)* 69+  0, 


(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  5+132, (2**17)*0+(2**8)*  8+ 79, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 15+106, (2**17)*0+(2**8)* 15+ 69, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 21+ 16, (2**17)*0+(2**8)* 26+145, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 37+142, (2**17)*0+(2**8)* 39+ 77, (2**17)*0+(2**8)* 71+150, (2**17)*1+(2**8)* 73+107, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  7+ 34, (2**17)*0+(2**8)* 12+  5, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 19+ 31, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 29+148, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 37+151, (2**17)*0+(2**8)* 37+ 93, (2**17)*0+(2**8)* 51+ 11, (2**17)*0+(2**8)* 60+ 79, (2**17)*0+(2**8)* 61+ 77, (2**17)*1+(2**8)* 67+  4, 
(2**17)*0+(2**8)*  3+132, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  9+141, (2**17)*0+(2**8)* 11+  7, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 21+155, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 40+ 53, (2**17)*0+(2**8)* 53+120, (2**17)*0+(2**8)* 54+ 91, (2**17)*0+(2**8)* 60+104, (2**17)*0+(2**8)* 68+ 66, (2**17)*1+(2**8)* 70+109, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  0+ 31, (2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 12+140, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 26+167, (2**17)*0+(2**8)* 27+ 27, (2**17)*0+(2**8)* 30+ 30, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 35+ 10, (2**17)*0+(2**8)* 55+  6, (2**17)*1+(2**8)* 57+ 99, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)*  4+ 13, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 10+ 60, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 17+ 33, (2**17)*0+(2**8)* 19+139, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 25+ 61, (2**17)*0+(2**8)* 28+ 14, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 33+  4, (2**17)*0+(2**8)* 36+165, (2**17)*0+(2**8)* 37+ 57, (2**17)*0+(2**8)* 37+ 45, (2**17)*0+(2**8)* 37+157, (2**17)*1+(2**8)* 43+147, 
(2**17)*0+(2**8)*  0+175, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  9+106, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 35+ 40, (2**17)*0+(2**8)* 37+ 21, (2**17)*0+(2**8)* 41+ 36, (2**17)*0+(2**8)* 48+151, (2**17)*0+(2**8)* 50+ 78, (2**17)*0+(2**8)* 50+ 99, (2**17)*0+(2**8)* 59+ 70, (2**17)*0+(2**8)* 59+ 79, (2**17)*1+(2**8)* 66+118, 
(2**17)*0+(2**8)*  0+ 79, (2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)*  1+120, (2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)* 10+ 10, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 20+145, (2**17)*0+(2**8)* 24+ 92, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 31+ 52, (2**17)*0+(2**8)* 32+124, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 39+ 26, (2**17)*0+(2**8)* 43+143, (2**17)*0+(2**8)* 55+ 61, (2**17)*1+(2**8)* 64+ 80, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 14+ 48, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 28+ 31, (2**17)*0+(2**8)* 34+ 59, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 37+ 35, (2**17)*0+(2**8)* 38+153, (2**17)*0+(2**8)* 42+149, (2**17)*0+(2**8)* 45+  9, (2**17)*0+(2**8)* 53+177, (2**17)*0+(2**8)* 62+157, (2**17)*1+(2**8)* 69+ 77, 
(2**17)*0+(2**8)*  0+141, (2**17)*0+(2**8)*  2+ 76, (2**17)*0+(2**8)* 34+149, (2**17)*0+(2**8)* 36+106, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 42+132, (2**17)*0+(2**8)* 45+ 79, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 52+106, (2**17)*0+(2**8)* 52+ 69, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 58+ 16, (2**17)*0+(2**8)* 63+145, (2**17)*1+(2**8)* 66+  0, 
(2**17)*0+(2**8)*  0+150, (2**17)*0+(2**8)*  0+ 92, (2**17)*0+(2**8)* 14+ 10, (2**17)*0+(2**8)* 23+ 78, (2**17)*0+(2**8)* 24+ 76, (2**17)*0+(2**8)* 30+  3, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 44+ 34, (2**17)*0+(2**8)* 49+  5, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 56+ 31, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 66+148, (2**17)*1+(2**8)* 67+  0, 
(2**17)*0+(2**8)*  3+ 52, (2**17)*0+(2**8)* 16+119, (2**17)*0+(2**8)* 17+ 90, (2**17)*0+(2**8)* 23+103, (2**17)*0+(2**8)* 31+ 65, (2**17)*0+(2**8)* 33+108, (2**17)*0+(2**8)* 40+132, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 46+141, (2**17)*0+(2**8)* 48+  7, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 58+155, (2**17)*0+(2**8)* 60+  0, (2**17)*1+(2**8)* 68+  0, 
(2**17)*0+(2**8)* 18+  5, (2**17)*0+(2**8)* 20+ 98, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 37+ 31, (2**17)*0+(2**8)* 44+ 51, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 49+140, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 63+167, (2**17)*0+(2**8)* 64+ 27, (2**17)*0+(2**8)* 67+ 30, (2**17)*0+(2**8)* 69+  0, (2**17)*1+(2**8)* 72+ 10, 
(2**17)*0+(2**8)*  0+ 56, (2**17)*0+(2**8)*  0+ 44, (2**17)*0+(2**8)*  0+156, (2**17)*0+(2**8)*  6+146, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 41+ 13, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 47+ 60, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 54+ 33, (2**17)*0+(2**8)* 56+139, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 62+ 61, (2**17)*0+(2**8)* 65+ 14, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 70+  4, (2**17)*1+(2**8)* 73+165, 
(2**17)*0+(2**8)*  0+ 20, (2**17)*0+(2**8)*  4+ 35, (2**17)*0+(2**8)* 11+150, (2**17)*0+(2**8)* 13+ 77, (2**17)*0+(2**8)* 13+ 98, (2**17)*0+(2**8)* 22+ 69, (2**17)*0+(2**8)* 22+ 78, (2**17)*0+(2**8)* 29+117, (2**17)*0+(2**8)* 37+175, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 46+106, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 71+  0, (2**17)*1+(2**8)* 72+ 40, 
(2**17)*0+(2**8)*  2+ 25, (2**17)*0+(2**8)*  6+142, (2**17)*0+(2**8)* 18+ 60, (2**17)*0+(2**8)* 27+ 79, (2**17)*0+(2**8)* 37+ 79, (2**17)*0+(2**8)* 37+106, (2**17)*0+(2**8)* 38+120, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 47+ 10, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 57+145, (2**17)*0+(2**8)* 61+ 92, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 68+ 52, (2**17)*0+(2**8)* 69+124, (2**17)*1+(2**8)* 72+  0, 
(2**17)*0+(2**8)*  0+ 34, (2**17)*0+(2**8)*  1+152, (2**17)*0+(2**8)*  5+148, (2**17)*0+(2**8)*  8+  8, (2**17)*0+(2**8)* 16+176, (2**17)*0+(2**8)* 25+156, (2**17)*0+(2**8)* 32+ 76, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 51+ 48, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 65+ 31, (2**17)*0+(2**8)* 71+ 59, (2**17)*1+(2**8)* 73+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  1+145, (2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  8+ 21, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 13+150, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 23+ 96, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 28+119, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 30+ 63, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 35+100, (2**17)*0+(2**8)* 40+ 81, (2**17)*0+(2**8)* 44+ 61, (2**17)*0+(2**8)* 48+120, (2**17)*0+(2**8)* 53+ 84, (2**17)*0+(2**8)* 56+116, (2**17)*0+(2**8)* 59+150, (2**17)*0+(2**8)* 60+ 39, (2**17)*0+(2**8)* 66+102, (2**17)*0+(2**8)* 74+116, (2**17)*1+(2**8)* 78+152, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)*  2+174, (2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  7+ 15, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 15+170, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 21+ 15, (2**17)*0+(2**8)* 24+145, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 27+126, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 31+ 42, (2**17)*0+(2**8)* 35+ 63, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 43+ 81, (2**17)*0+(2**8)* 43+157, (2**17)*0+(2**8)* 45+ 93, (2**17)*0+(2**8)* 52+137, (2**17)*0+(2**8)* 54+150, (2**17)*0+(2**8)* 55+101, (2**17)*0+(2**8)* 69+125, (2**17)*0+(2**8)* 74+ 56, (2**17)*1+(2**8)* 78+ 51, 
(2**17)*0+(2**8)*  0+ 71, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  4+ 48, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  9+ 69, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 14+ 50, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 22+ 20, (2**17)*0+(2**8)* 25+172, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 29+147, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 33+ 39, (2**17)*0+(2**8)* 36+ 73, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 39+117, (2**17)*0+(2**8)* 41+134, (2**17)*0+(2**8)* 46+ 78, (2**17)*0+(2**8)* 50+ 43, (2**17)*0+(2**8)* 56+ 10, (2**17)*0+(2**8)* 57+ 66, (2**17)*0+(2**8)* 61+ 37, (2**17)*1+(2**8)* 73+ 58, 
(2**17)*0+(2**8)*  1+ 87, (2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  4+ 92, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 17+140, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 18+145, (2**17)*0+(2**8)* 22+132, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 40+156, (2**17)*0+(2**8)* 45+158, (2**17)*0+(2**8)* 47+ 61, (2**17)*0+(2**8)* 50+ 49, (2**17)*0+(2**8)* 51+ 83, (2**17)*0+(2**8)* 63+ 32, (2**17)*0+(2**8)* 65+110, (2**17)*0+(2**8)* 66+143, (2**17)*0+(2**8)* 70+ 51, (2**17)*0+(2**8)* 72+ 90, (2**17)*0+(2**8)* 76+137, (2**17)*1+(2**8)* 77+133, 
(2**17)*0+(2**8)*  2+118, (2**17)*0+(2**8)*  3+ 29, (2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)*  6+137, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)*  9+148, (2**17)*0+(2**8)* 11+112, (2**17)*0+(2**8)* 12+ 87, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 18+ 62, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 27+156, (2**17)*0+(2**8)* 28+ 54, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 31+170, (2**17)*0+(2**8)* 32+ 28, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 39+110, (2**17)*0+(2**8)* 42+113, (2**17)*0+(2**8)* 59+ 43, (2**17)*0+(2**8)* 60+ 81, (2**17)*0+(2**8)* 64+104, (2**17)*1+(2**8)* 77+ 33, 
(2**17)*0+(2**8)*  0+ 80, (2**17)*0+(2**8)*  4+ 60, (2**17)*0+(2**8)*  8+119, (2**17)*0+(2**8)* 13+ 83, (2**17)*0+(2**8)* 16+115, (2**17)*0+(2**8)* 19+149, (2**17)*0+(2**8)* 20+ 38, (2**17)*0+(2**8)* 26+101, (2**17)*0+(2**8)* 34+115, (2**17)*0+(2**8)* 38+151, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 41+145, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 48+ 21, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 53+150, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 63+ 96, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 68+119, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 70+ 63, (2**17)*0+(2**8)* 75+  0, (2**17)*1+(2**8)* 75+100, 
(2**17)*0+(2**8)*  3+ 80, (2**17)*0+(2**8)*  3+156, (2**17)*0+(2**8)*  5+ 92, (2**17)*0+(2**8)* 12+136, (2**17)*0+(2**8)* 14+149, (2**17)*0+(2**8)* 15+100, (2**17)*0+(2**8)* 29+124, (2**17)*0+(2**8)* 34+ 55, (2**17)*0+(2**8)* 38+ 50, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 42+174, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 47+ 15, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 55+170, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 61+ 15, (2**17)*0+(2**8)* 64+145, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 67+126, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 71+ 42, (2**17)*0+(2**8)* 75+ 63, (2**17)*1+(2**8)* 76+  0, 
(2**17)*0+(2**8)*  1+133, (2**17)*0+(2**8)*  6+ 77, (2**17)*0+(2**8)* 10+ 42, (2**17)*0+(2**8)* 16+  9, (2**17)*0+(2**8)* 17+ 65, (2**17)*0+(2**8)* 21+ 36, (2**17)*0+(2**8)* 33+ 57, (2**17)*0+(2**8)* 40+ 71, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 44+ 48, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 49+ 69, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 54+ 50, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 62+ 20, (2**17)*0+(2**8)* 65+172, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 69+147, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 73+ 39, (2**17)*0+(2**8)* 76+ 73, (2**17)*0+(2**8)* 77+  0, (2**17)*1+(2**8)* 79+117, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)*  5+157, (2**17)*0+(2**8)*  7+ 60, (2**17)*0+(2**8)* 10+ 48, (2**17)*0+(2**8)* 11+ 82, (2**17)*0+(2**8)* 23+ 31, (2**17)*0+(2**8)* 25+109, (2**17)*0+(2**8)* 26+142, (2**17)*0+(2**8)* 30+ 50, (2**17)*0+(2**8)* 32+ 89, (2**17)*0+(2**8)* 36+136, (2**17)*0+(2**8)* 37+132, (2**17)*0+(2**8)* 41+ 87, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 44+ 92, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 57+140, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 58+145, (2**17)*0+(2**8)* 62+132, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 73+  0, (2**17)*1+(2**8)* 78+  0, 
(2**17)*0+(2**8)*  2+112, (2**17)*0+(2**8)* 19+ 42, (2**17)*0+(2**8)* 20+ 80, (2**17)*0+(2**8)* 24+103, (2**17)*0+(2**8)* 37+ 32, (2**17)*0+(2**8)* 42+118, (2**17)*0+(2**8)* 43+ 29, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 46+137, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 49+148, (2**17)*0+(2**8)* 51+112, (2**17)*0+(2**8)* 52+ 87, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 58+ 62, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 67+156, (2**17)*0+(2**8)* 68+ 54, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 71+170, (2**17)*0+(2**8)* 72+ 28, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 79+  0, (2**17)*1+(2**8)* 79+110, 


(2**17)*0+(2**8)*  0+  2, (2**17)*1+(2**8)* 72+ 35, 
(2**17)*0+(2**8)* 73+134, (2**17)*1+(2**8)* 89+122, 
(2**17)*0+(2**8)*  6+  7, (2**17)*1+(2**8)* 14+ 10, 
(2**17)*0+(2**8)* 13+166, (2**17)*1+(2**8)* 65+163, 
(2**17)*0+(2**8)* 46+ 62, (2**17)*1+(2**8)* 56+178, 
(2**17)*0+(2**8)* 49+101, (2**17)*1+(2**8)* 70+163, 
(2**17)*0+(2**8)* 50+ 52, (2**17)*1+(2**8)* 50+ 95, 
(2**17)*0+(2**8)* 55+ 51, (2**17)*1+(2**8)* 57+156, 
(2**17)*0+(2**8)* 24+143, (2**17)*1+(2**8)* 35+113, 
(2**17)*0+(2**8)* 62+ 24, (2**17)*1+(2**8)* 86+110, 
(2**17)*0+(2**8)*  9+156, (2**17)*1+(2**8)* 55+ 32, 
(2**17)*0+(2**8)* 12+ 31, (2**17)*1+(2**8)* 47+ 49, 
(2**17)*0+(2**8)* 15+ 82, (2**17)*1+(2**8)* 53+112, 
(2**17)*0+(2**8)* 59+119, (2**17)*1+(2**8)* 87+122, 
(2**17)*0+(2**8)* 11+ 72, (2**17)*1+(2**8)* 29+ 27, 
(2**17)*0+(2**8)*  2+112, (2**17)*1+(2**8)* 45+ 69, 
(2**17)*0+(2**8)*  0+ 23, (2**17)*1+(2**8)*  7+164, 
(2**17)*0+(2**8)*  8+162, (2**17)*1+(2**8)* 12+ 46, 
(2**17)*0+(2**8)*  9+103, (2**17)*1+(2**8)* 40+ 63, 
(2**17)*0+(2**8)* 53+155, (2**17)*1+(2**8)* 57+ 98, 
(2**17)*0+(2**8)* 11+163, (2**17)*1+(2**8)* 30+ 48, 
(2**17)*0+(2**8)* 59+102, (2**17)*1+(2**8)* 68+ 90, 
(2**17)*0+(2**8)* 46+ 93, (2**17)*1+(2**8)* 80+137, 
(2**17)*0+(2**8)* 10+ 96, (2**17)*1+(2**8)* 36+ 28, 
(2**17)*0+(2**8)*  8+107, (2**17)*1+(2**8)* 51+167, 
(2**17)*0+(2**8)*  5+ 83, (2**17)*1+(2**8)* 58+139, 
(2**17)*0+(2**8)* 62+130, (2**17)*1+(2**8)* 79+ 91, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*1+(2**8)* 49+107, 
(2**17)*0+(2**8)*  7+149, (2**17)*1+(2**8)* 59+144, 
(2**17)*0+(2**8)* 45+156, (2**17)*1+(2**8)* 47+ 54, 
(2**17)*0+(2**8)*  6+156, (2**17)*1+(2**8)* 75+ 63, 
(2**17)*0+(2**8)*  4+ 37, (2**17)*1+(2**8)*  5+121, 
(2**17)*0+(2**8)* 36+ 90, (2**17)*1+(2**8)* 69+115, 
(2**17)*0+(2**8)* 11+ 90, (2**17)*1+(2**8)* 70+132, 
(2**17)*0+(2**8)*  1+137, (2**17)*1+(2**8)*  8+ 80, 
(2**17)*0+(2**8)* 55+115, (2**17)*1+(2**8)* 85+ 35, 
(2**17)*0+(2**8)* 49+150, (2**17)*1+(2**8)* 51+ 86, 
(2**17)*0+(2**8)* 46+ 77, (2**17)*1+(2**8)* 54+127, 
(2**17)*0+(2**8)*  3+148, (2**17)*1+(2**8)* 27+ 81, 
(2**17)*0+(2**8)* 19+ 53, (2**17)*1+(2**8)* 54+ 17, 
(2**17)*0+(2**8)*  5+150, (2**17)*1+(2**8)* 78+ 33, 
(2**17)*0+(2**8)* 13+ 50, (2**17)*1+(2**8)* 58+ 87, 
(2**17)*0+(2**8)*  0+ 88, (2**17)*1+(2**8)* 61+ 72, 
(2**17)*0+(2**8)* 66+ 32, (2**17)*1+(2**8)* 82+  2, 
(2**17)*0+(2**8)*  9+ 14, (2**17)*1+(2**8)* 47+ 43, 
(2**17)*0+(2**8)*  5+ 68, (2**17)*1+(2**8)* 53+ 78, 
(2**17)*0+(2**8)* 12+101, (2**17)*1+(2**8)* 51+ 19, 
(2**17)*0+(2**8)*  7+ 51, (2**17)*1+(2**8)* 64+180, 
(2**17)*0+(2**8)*  6+ 38, (2**17)*1+(2**8)* 11+ 63, 
(2**17)*0+(2**8)* 13+172, (2**17)*1+(2**8)* 56+ 72, 
(2**17)*0+(2**8)*  4+ 50, (2**17)*1+(2**8)* 31+ 83, 
(2**17)*0+(2**8)*  7+139, (2**17)*1+(2**8)* 58+ 12, 
(2**17)*0+(2**8)*  4+155, (2**17)*1+(2**8)*  8+ 42, 
(2**17)*0+(2**8)* 13+131, (2**17)*1+(2**8)* 45+134, 
(2**17)*0+(2**8)* 11+ 56, (2**17)*1+(2**8)* 68+ 76, 
(2**17)*0+(2**8)*  2+115, (2**17)*1+(2**8)* 67+ 89, 
(2**17)*0+(2**8)* 37+100, (2**17)*1+(2**8)* 67+107, 
(2**17)*0+(2**8)* 51+ 33, (2**17)*1+(2**8)* 54+141, 
(2**17)*0+(2**8)*  0+ 67, (2**17)*1+(2**8)* 38+116, 
(2**17)*0+(2**8)*  2+143, (2**17)*1+(2**8)* 48+ 23, 
(2**17)*0+(2**8)*  0+  4, (2**17)*1+(2**8)*  7+ 44, 
(2**17)*0+(2**8)* 39+  8, (2**17)*1+(2**8)* 56+ 16, 
(2**17)*0+(2**8)* 46+158, (2**17)*1+(2**8)* 60+ 31, 
(2**17)*0+(2**8)* 41+ 64, (2**17)*1+(2**8)* 59+159, 
(2**17)*0+(2**8)*  3+150, (2**17)*1+(2**8)* 13+ 33, 
(2**17)*0+(2**8)* 51+ 59, (2**17)*1+(2**8)* 56+160, 
(2**17)*0+(2**8)* 33+175, (2**17)*1+(2**8)* 58+ 22, 
(2**17)*0+(2**8)*  8+ 24, (2**17)*1+(2**8)* 57+ 68, 
(2**17)*0+(2**8)* 56+ 18, (2**17)*1+(2**8)* 83+ 45, 
(2**17)*0+(2**8)*  9+ 21, (2**17)*1+(2**8)* 35+  3, 
(2**17)*0+(2**8)*  8+104, (2**17)*1+(2**8)* 38+ 80, 
(2**17)*0+(2**8)* 26+ 26, (2**17)*1+(2**8)* 47+107, 
(2**17)*0+(2**8)* 49+ 30, (2**17)*1+(2**8)* 79+ 56, 
(2**17)*0+(2**8)*  5+145, (2**17)*1+(2**8)* 52+ 39, 
(2**17)*0+(2**8)*  2+ 69, (2**17)*1+(2**8)*  4+ 49, 
(2**17)*0+(2**8)* 10+145, (2**17)*1+(2**8)* 54+101, 
(2**17)*0+(2**8)* 12+172, (2**17)*1+(2**8)* 84+ 67, 
(2**17)*0+(2**8)*  5+ 46, (2**17)*1+(2**8)* 57+110, 
(2**17)*0+(2**8)* 59+143, (2**17)*1+(2**8)* 71+ 56, 
(2**17)*0+(2**8)* 11+ 70, (2**17)*1+(2**8)* 39+  4, 
(2**17)*0+(2**8)*  4+170, (2**17)*1+(2**8)*  6+169, 
(2**17)*0+(2**8)* 11+109, (2**17)*1+(2**8)* 17+124, 
(2**17)*0+(2**8)* 18+110, (2**17)*1+(2**8)* 77+ 37, 
(2**17)*0+(2**8)* 48+ 58, (2**17)*1+(2**8)* 50+165, 
(2**17)*0+(2**8)* 46+ 61, (2**17)*1+(2**8)* 76+ 88, 
(2**17)*0+(2**8)*  8+  3, (2**17)*1+(2**8)* 77+165, 
(2**17)*0+(2**8)*  4+ 72, (2**17)*1+(2**8)*  8+ 95, 
(2**17)*0+(2**8)* 24+ 30, (2**17)*1+(2**8)* 52+122, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*1+(2**8)* 47+ 83, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*1+(2**8)* 57+ 62, 
(2**17)*0+(2**8)* 53+ 25, (2**17)*1+(2**8)* 57+ 35, 
(2**17)*0+(2**8)*  1+129, (2**17)*1+(2**8)* 73+ 44, 
(2**17)*0+(2**8)* 29+147, (2**17)*1+(2**8)* 37+ 17, 
(2**17)*0+(2**8)* 18+109, (2**17)*1+(2**8)* 87+171, 
(2**17)*0+(2**8)* 12+119, (2**17)*1+(2**8)* 48+115, 
(2**17)*0+(2**8)* 18+114, (2**17)*1+(2**8)* 86+ 91, 
(2**17)*0+(2**8)* 12+131, (2**17)*1+(2**8)* 60+ 90, 
(2**17)*0+(2**8)* 14+ 77, (2**17)*1+(2**8)* 66+123, 
(2**17)*0+(2**8)*  7+172, (2**17)*1+(2**8)* 19+ 34, 
(2**17)*0+(2**8)*  9+132, (2**17)*1+(2**8)* 47+ 52, 
(2**17)*0+(2**8)* 10+ 12, (2**17)*1+(2**8)* 48+ 84, 
(2**17)*0+(2**8)*  7+ 13, (2**17)*1+(2**8)* 31+ 41, 
(2**17)*0+(2**8)* 44+ 76, (2**17)*1+(2**8)* 58+ 27, 
(2**17)*0+(2**8)* 46+ 64, (2**17)*1+(2**8)* 55+118, 
(2**17)*0+(2**8)* 45+107, (2**17)*1+(2**8)* 50+148, 
(2**17)*0+(2**8)* 27+ 20, (2**17)*1+(2**8)* 40+143, 
(2**17)*0+(2**8)* 55+127, (2**17)*1+(2**8)* 74+125, 
(2**17)*0+(2**8)* 10+ 32, (2**17)*1+(2**8)* 59+153, 
(2**17)*0+(2**8)*  0+174, (2**17)*1+(2**8)* 51+168, 
(2**17)*0+(2**8)*  4+ 91, (2**17)*1+(2**8)* 73+122, 
(2**17)*0+(2**8)* 14+ 98, (2**17)*1+(2**8)* 89+173, 
(2**17)*0+(2**8)* 10+  4, (2**17)*1+(2**8)* 51+ 72, 
(2**17)*0+(2**8)* 68+ 15, (2**17)*1+(2**8)* 88+137, 
(2**17)*0+(2**8)*  6+ 56, (2**17)*1+(2**8)* 54+ 26, 
(2**17)*0+(2**8)*  3+ 82, (2**17)*1+(2**8)*  3+ 62, 
(2**17)*0+(2**8)*  9+ 40, (2**17)*1+(2**8)* 20+ 15, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*1+(2**8)* 77+128, 
(2**17)*0+(2**8)* 46+ 78, (2**17)*1+(2**8)* 58+ 58, 
(2**17)*0+(2**8)*  1+ 62, (2**17)*1+(2**8)* 55+ 47, 
(2**17)*0+(2**8)* 14+  5, (2**17)*1+(2**8)* 47+  7, 
(2**17)*0+(2**8)* 21+127, (2**17)*1+(2**8)* 88+ 68, 
(2**17)*0+(2**8)* 55+ 62, (2**17)*1+(2**8)* 71+169, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*1+(2**8)* 34+168, 
(2**17)*0+(2**8)* 43+ 75, (2**17)*1+(2**8)* 61+ 37, 
(2**17)*0+(2**8)*  7+119, (2**17)*1+(2**8)* 87+115, 
(2**17)*0+(2**8)* 22+ 83, (2**17)*1+(2**8)* 59+101, 
(2**17)*0+(2**8)*  4+121, (2**17)*1+(2**8)* 65+141, 
(2**17)*0+(2**8)* 61+103, (2**17)*1+(2**8)* 75+111, 
(2**17)*0+(2**8)* 50+129, (2**17)*1+(2**8)* 58+ 99, 
(2**17)*0+(2**8)* 25+ 79, (2**17)*1+(2**8)* 59+174, 
(2**17)*0+(2**8)*  7+  5, (2**17)*1+(2**8)* 78+ 52, 
(2**17)*0+(2**8)*  5+ 36, (2**17)*1+(2**8)* 48+ 34, 
(2**17)*0+(2**8)*  3+ 88, (2**17)*1+(2**8)*  9+ 81, 
(2**17)*0+(2**8)*  1+ 28, (2**17)*1+(2**8)*  7+ 25, 
(2**17)*0+(2**8)*  2+148, (2**17)*1+(2**8)* 36+ 49, 
(2**17)*0+(2**8)* 27+ 34, (2**17)*1+(2**8)* 45+  2, 
(2**17)*0+(2**8)* 28+133, (2**17)*1+(2**8)* 44+121, 
(2**17)*0+(2**8)* 51+  7, (2**17)*1+(2**8)* 59+ 10, 
(2**17)*0+(2**8)* 20+162, (2**17)*1+(2**8)* 58+166, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*1+(2**8)* 11+177, 
(2**17)*0+(2**8)*  4+100, (2**17)*1+(2**8)* 25+162, 
(2**17)*0+(2**8)*  5+ 51, (2**17)*1+(2**8)*  5+ 94, 
(2**17)*0+(2**8)* 10+ 50, (2**17)*1+(2**8)* 12+155, 
(2**17)*0+(2**8)* 69+143, (2**17)*1+(2**8)* 80+113, 
(2**17)*0+(2**8)* 17+ 23, (2**17)*1+(2**8)* 41+109, 
(2**17)*0+(2**8)* 10+ 31, (2**17)*1+(2**8)* 54+156, 
(2**17)*0+(2**8)*  2+ 48, (2**17)*1+(2**8)* 57+ 31, 
(2**17)*0+(2**8)*  8+111, (2**17)*1+(2**8)* 60+ 82, 
(2**17)*0+(2**8)* 14+118, (2**17)*1+(2**8)* 42+121, 
(2**17)*0+(2**8)* 56+ 72, (2**17)*1+(2**8)* 74+ 27, 
(2**17)*0+(2**8)*  0+ 68, (2**17)*1+(2**8)* 47+112, 
(2**17)*0+(2**8)* 45+ 23, (2**17)*1+(2**8)* 52+164, 
(2**17)*0+(2**8)* 53+162, (2**17)*1+(2**8)* 57+ 46, 
(2**17)*0+(2**8)* 54+103, (2**17)*1+(2**8)* 85+ 63, 
(2**17)*0+(2**8)*  8+154, (2**17)*1+(2**8)* 12+ 97, 
(2**17)*0+(2**8)* 56+163, (2**17)*1+(2**8)* 75+ 48, 
(2**17)*0+(2**8)* 14+101, (2**17)*1+(2**8)* 23+ 89, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*1+(2**8)* 35+136, 
(2**17)*0+(2**8)* 55+ 96, (2**17)*1+(2**8)* 81+ 28, 
(2**17)*0+(2**8)*  6+166, (2**17)*1+(2**8)* 53+107, 
(2**17)*0+(2**8)* 13+138, (2**17)*1+(2**8)* 50+ 83, 
(2**17)*0+(2**8)* 17+129, (2**17)*1+(2**8)* 34+ 90, 
(2**17)*0+(2**8)*  4+106, (2**17)*1+(2**8)* 48+ 33, 
(2**17)*0+(2**8)* 14+143, (2**17)*1+(2**8)* 52+149, 
(2**17)*0+(2**8)*  0+155, (2**17)*1+(2**8)*  2+ 53, 
(2**17)*0+(2**8)* 30+ 62, (2**17)*1+(2**8)* 51+156, 
(2**17)*0+(2**8)* 49+ 37, (2**17)*1+(2**8)* 50+121, 
(2**17)*0+(2**8)* 24+114, (2**17)*1+(2**8)* 81+ 90, 
(2**17)*0+(2**8)* 25+131, (2**17)*1+(2**8)* 56+ 90, 
(2**17)*0+(2**8)* 46+137, (2**17)*1+(2**8)* 53+ 80, 
(2**17)*0+(2**8)* 10+114, (2**17)*1+(2**8)* 40+ 34, 
(2**17)*0+(2**8)*  4+149, (2**17)*1+(2**8)*  6+ 85, 
(2**17)*0+(2**8)*  1+ 76, (2**17)*1+(2**8)*  9+126, 
(2**17)*0+(2**8)* 48+148, (2**17)*1+(2**8)* 72+ 81, 
(2**17)*0+(2**8)*  9+ 16, (2**17)*1+(2**8)* 64+ 53, 
(2**17)*0+(2**8)* 33+ 32, (2**17)*1+(2**8)* 50+150, 
(2**17)*0+(2**8)* 13+ 86, (2**17)*1+(2**8)* 58+ 50, 
(2**17)*0+(2**8)* 16+ 71, (2**17)*1+(2**8)* 45+ 88, 
(2**17)*0+(2**8)* 21+ 31, (2**17)*1+(2**8)* 37+  1, 
(2**17)*0+(2**8)*  2+ 42, (2**17)*1+(2**8)* 54+ 14, 
(2**17)*0+(2**8)*  8+ 77, (2**17)*1+(2**8)* 50+ 68, 
(2**17)*0+(2**8)*  6+ 18, (2**17)*1+(2**8)* 57+101, 
(2**17)*0+(2**8)* 19+179, (2**17)*1+(2**8)* 52+ 51, 
(2**17)*0+(2**8)* 51+ 38, (2**17)*1+(2**8)* 56+ 63, 
(2**17)*0+(2**8)* 11+ 71, (2**17)*1+(2**8)* 58+172, 
(2**17)*0+(2**8)* 49+ 50, (2**17)*1+(2**8)* 76+ 83, 
(2**17)*0+(2**8)* 13+ 11, (2**17)*1+(2**8)* 52+139, 
(2**17)*0+(2**8)* 49+155, (2**17)*1+(2**8)* 53+ 42, 
(2**17)*0+(2**8)*  0+133, (2**17)*1+(2**8)* 58+131, 
(2**17)*0+(2**8)* 23+ 75, (2**17)*1+(2**8)* 56+ 56, 
(2**17)*0+(2**8)* 22+ 88, (2**17)*1+(2**8)* 47+115, 
(2**17)*0+(2**8)* 22+106, (2**17)*1+(2**8)* 82+100, 
(2**17)*0+(2**8)*  6+ 32, (2**17)*1+(2**8)*  9+140, 
(2**17)*0+(2**8)* 45+ 67, (2**17)*1+(2**8)* 83+116, 
(2**17)*0+(2**8)*  3+ 22, (2**17)*1+(2**8)* 47+143, 
(2**17)*0+(2**8)* 45+  4, (2**17)*1+(2**8)* 52+ 44, 
(2**17)*0+(2**8)* 11+ 15, (2**17)*1+(2**8)* 84+  8, 
(2**17)*0+(2**8)*  1+157, (2**17)*1+(2**8)* 15+ 30, 
(2**17)*0+(2**8)* 14+158, (2**17)*1+(2**8)* 86+ 64, 
(2**17)*0+(2**8)* 48+150, (2**17)*1+(2**8)* 58+ 33, 
(2**17)*0+(2**8)*  6+ 58, (2**17)*1+(2**8)* 11+159, 
(2**17)*0+(2**8)* 13+ 21, (2**17)*1+(2**8)* 78+175, 
(2**17)*0+(2**8)* 12+ 67, (2**17)*1+(2**8)* 53+ 24, 
(2**17)*0+(2**8)* 11+ 17, (2**17)*1+(2**8)* 38+ 44, 
(2**17)*0+(2**8)* 54+ 21, (2**17)*1+(2**8)* 80+  3, 
(2**17)*0+(2**8)* 53+104, (2**17)*1+(2**8)* 83+ 80, 
(2**17)*0+(2**8)*  2+106, (2**17)*1+(2**8)* 71+ 26, 
(2**17)*0+(2**8)*  4+ 29, (2**17)*1+(2**8)* 34+ 55, 
(2**17)*0+(2**8)*  7+ 38, (2**17)*1+(2**8)* 50+145, 
(2**17)*0+(2**8)* 47+ 69, (2**17)*1+(2**8)* 49+ 49, 
(2**17)*0+(2**8)*  9+100, (2**17)*1+(2**8)* 55+145, 
(2**17)*0+(2**8)* 39+ 66, (2**17)*1+(2**8)* 57+172, 
(2**17)*0+(2**8)* 12+109, (2**17)*1+(2**8)* 50+ 46, 
(2**17)*0+(2**8)* 14+142, (2**17)*1+(2**8)* 26+ 55, 
(2**17)*0+(2**8)* 56+ 70, (2**17)*1+(2**8)* 84+  4, 
(2**17)*0+(2**8)* 49+170, (2**17)*1+(2**8)* 51+169, 
(2**17)*0+(2**8)* 56+109, (2**17)*1+(2**8)* 62+124, 
(2**17)*0+(2**8)* 32+ 36, (2**17)*1+(2**8)* 63+110, 
(2**17)*0+(2**8)*  3+ 57, (2**17)*1+(2**8)*  5+164, 
(2**17)*0+(2**8)*  1+ 60, (2**17)*1+(2**8)* 31+ 87, 
(2**17)*0+(2**8)* 32+164, (2**17)*1+(2**8)* 53+  3, 
(2**17)*0+(2**8)* 49+ 72, (2**17)*1+(2**8)* 53+ 95, 
(2**17)*0+(2**8)*  7+121, (2**17)*1+(2**8)* 69+ 30, 
(2**17)*0+(2**8)*  2+ 82, (2**17)*1+(2**8)* 46+ 92, 
(2**17)*0+(2**8)* 12+ 61, (2**17)*1+(2**8)* 45+ 77, 
(2**17)*0+(2**8)*  8+ 24, (2**17)*1+(2**8)* 12+ 34, 
(2**17)*0+(2**8)* 28+ 43, (2**17)*1+(2**8)* 46+129, 
(2**17)*0+(2**8)* 74+147, (2**17)*1+(2**8)* 82+ 17, 
(2**17)*0+(2**8)* 42+170, (2**17)*1+(2**8)* 63+109, 
(2**17)*0+(2**8)*  3+114, (2**17)*1+(2**8)* 57+119, 
(2**17)*0+(2**8)* 41+ 90, (2**17)*1+(2**8)* 63+114, 
(2**17)*0+(2**8)* 15+ 89, (2**17)*1+(2**8)* 57+131, 
(2**17)*0+(2**8)* 21+122, (2**17)*1+(2**8)* 59+ 77, 
(2**17)*0+(2**8)* 52+172, (2**17)*1+(2**8)* 64+ 34, 
(2**17)*0+(2**8)*  2+ 51, (2**17)*1+(2**8)* 54+132, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*1+(2**8)* 55+ 12, 
(2**17)*0+(2**8)* 52+ 13, (2**17)*1+(2**8)* 76+ 41, 
(2**17)*0+(2**8)* 13+ 26, (2**17)*1+(2**8)* 89+ 76, 
(2**17)*0+(2**8)*  1+ 63, (2**17)*1+(2**8)* 10+117, 
(2**17)*0+(2**8)*  0+106, (2**17)*1+(2**8)*  5+147, 
(2**17)*0+(2**8)* 72+ 20, (2**17)*1+(2**8)* 85+143, 
(2**17)*0+(2**8)* 10+126, (2**17)*1+(2**8)* 29+124, 
(2**17)*0+(2**8)* 14+152, (2**17)*1+(2**8)* 55+ 32, 
(2**17)*0+(2**8)*  6+167, (2**17)*1+(2**8)* 45+174, 
(2**17)*0+(2**8)* 28+121, (2**17)*1+(2**8)* 49+ 91, 
(2**17)*0+(2**8)* 44+172, (2**17)*1+(2**8)* 59+ 98, 
(2**17)*0+(2**8)*  6+ 71, (2**17)*1+(2**8)* 55+  4, 
(2**17)*0+(2**8)* 23+ 14, (2**17)*1+(2**8)* 43+136, 
(2**17)*0+(2**8)*  9+ 25, (2**17)*1+(2**8)* 51+ 56, 
(2**17)*0+(2**8)* 48+ 82, (2**17)*1+(2**8)* 48+ 62, 
(2**17)*0+(2**8)* 54+ 40, (2**17)*1+(2**8)* 65+ 15, 
(2**17)*0+(2**8)* 32+127, (2**17)*1+(2**8)* 45+ 87, 
(2**17)*0+(2**8)*  1+ 77, (2**17)*1+(2**8)* 13+ 57, 
(2**17)*0+(2**8)* 10+ 46, (2**17)*1+(2**8)* 46+ 62, 
(2**17)*0+(2**8)*  2+  6, (2**17)*1+(2**8)* 59+  5, 
(2**17)*0+(2**8)* 43+ 67, (2**17)*1+(2**8)* 66+127, 
(2**17)*0+(2**8)* 10+ 61, (2**17)*1+(2**8)* 26+168, 
(2**17)*0+(2**8)* 48+ 83, (2**17)*1+(2**8)* 79+168, 
(2**17)*0+(2**8)* 16+ 36, (2**17)*1+(2**8)* 88+ 75, 
(2**17)*0+(2**8)* 42+114, (2**17)*1+(2**8)* 52+119, 
(2**17)*0+(2**8)* 14+100, (2**17)*1+(2**8)* 67+ 83, 
(2**17)*0+(2**8)* 20+140, (2**17)*1+(2**8)* 49+121, 
(2**17)*0+(2**8)* 16+102, (2**17)*1+(2**8)* 30+110, 
(2**17)*0+(2**8)*  5+128, (2**17)*1+(2**8)* 13+ 98, 
(2**17)*0+(2**8)* 14+173, (2**17)*1+(2**8)* 70+ 79, 
(2**17)*0+(2**8)* 33+ 51, (2**17)*1+(2**8)* 52+  5, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*1+(2**8)* 50+ 36, 
(2**17)*0+(2**8)* 48+ 88, (2**17)*1+(2**8)* 54+ 81, 
(2**17)*0+(2**8)* 46+ 28, (2**17)*1+(2**8)* 52+ 25, 
(2**17)*0+(2**8)* 47+148, (2**17)*1+(2**8)* 81+ 49, 


(2**17)*0+(2**8)*  0+ 23, (2**17)*0+(2**8)*  0+ 88, (2**17)*1+(2**8)*104+157, 
(2**17)*0+(2**8)* 35+114, (2**17)*0+(2**8)* 46+ 92, (2**17)*1+(2**8)* 54+118, 
(2**17)*0+(2**8)* 27+142, (2**17)*0+(2**8)* 66+ 72, (2**17)*1+(2**8)* 76+122, 
(2**17)*0+(2**8)* 12+166, (2**17)*0+(2**8)* 61+ 62, (2**17)*1+(2**8)*106+105, 
(2**17)*0+(2**8)* 13+ 10, (2**17)*0+(2**8)* 70+178, (2**17)*1+(2**8)* 83+173, 
(2**17)*0+(2**8)* 17+ 43, (2**17)*0+(2**8)* 18+  8, (2**17)*1+(2**8)* 64+101, 
(2**17)*0+(2**8)* 65+ 52, (2**17)*0+(2**8)* 65+ 95, (2**17)*1+(2**8)* 75+132, 
(2**17)*0+(2**8)* 18+ 64, (2**17)*0+(2**8)* 69+ 51, (2**17)*1+(2**8)*107+ 34, 
(2**17)*0+(2**8)* 34+165, (2**17)*0+(2**8)* 81+ 73, (2**17)*1+(2**8)* 82+ 67, 
(2**17)*0+(2**8)* 16+ 27, (2**17)*0+(2**8)* 69+145, (2**17)*1+(2**8)* 83+114, 
(2**17)*0+(2**8)* 62+ 49, (2**17)*0+(2**8)* 79+ 89, (2**17)*1+(2**8)*105+132, 
(2**17)*0+(2**8)*  8+156, (2**17)*0+(2**8)* 16+ 54, (2**17)*1+(2**8)* 69+ 32, 
(2**17)*0+(2**8)* 74+ 76, (2**17)*0+(2**8)* 76+156, (2**17)*1+(2**8)*114+ 21, 
(2**17)*0+(2**8)*  0+ 67, (2**17)*0+(2**8)* 10+ 72, (2**17)*1+(2**8)* 11+ 31, 
(2**17)*0+(2**8)*  2+112, (2**17)*0+(2**8)* 60+ 69, (2**17)*1+(2**8)* 82+162, 
(2**17)*0+(2**8)*  7+164, (2**17)*0+(2**8)* 11+ 46, (2**17)*1+(2**8)*104+ 60, 
(2**17)*0+(2**8)* 17+  3, (2**17)*0+(2**8)* 52+  5, (2**17)*1+(2**8)* 57+ 33, 
(2**17)*0+(2**8)* 34+ 88, (2**17)*0+(2**8)* 73+119, (2**17)*1+(2**8)* 95+123, 
(2**17)*0+(2**8)*  8+103, (2**17)*0+(2**8)* 58+ 44, (2**17)*1+(2**8)* 67+131, 
(2**17)*0+(2**8)* 10+163, (2**17)*0+(2**8)* 82+119, (2**17)*1+(2**8)*106+106, 
(2**17)*0+(2**8)* 32+166, (2**17)*0+(2**8)* 70+ 49, (2**17)*1+(2**8)* 74+ 32, 
(2**17)*0+(2**8)* 16+119, (2**17)*0+(2**8)* 65+170, (2**17)*1+(2**8)* 71+ 98, 
(2**17)*0+(2**8)* 61+ 93, (2**17)*0+(2**8)* 67+ 81, (2**17)*1+(2**8)* 72+139, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*0+(2**8)* 29+ 74, (2**17)*1+(2**8)* 77+ 37, 
(2**17)*0+(2**8)*  9+ 96, (2**17)*0+(2**8)* 37+ 80, (2**17)*1+(2**8)*103+ 78, 
(2**17)*0+(2**8)* 15+ 79, (2**17)*0+(2**8)* 18+119, (2**17)*1+(2**8)* 66+ 19, 
(2**17)*0+(2**8)*  0+  2, (2**17)*0+(2**8)*  5+ 83, (2**17)*1+(2**8)*  8+127, 
(2**17)*0+(2**8)*  7+149, (2**17)*0+(2**8)* 55+ 17, (2**17)*1+(2**8)* 62+ 54, 
(2**17)*0+(2**8)* 17+ 48, (2**17)*0+(2**8)* 64+107, (2**17)*1+(2**8)*117+162, 
(2**17)*0+(2**8)* 41+107, (2**17)*0+(2**8)* 73+ 94, (2**17)*1+(2**8)* 80+118, 
(2**17)*0+(2**8)*  1+137, (2**17)*0+(2**8)*  6+169, (2**17)*1+(2**8)* 76+ 73, 
(2**17)*0+(2**8)* 64+150, (2**17)*0+(2**8)* 73+144, (2**17)*1+(2**8)*119+166, 
(2**17)*0+(2**8)*  5+121, (2**17)*0+(2**8)*  6+  7, (2**17)*1+(2**8)* 79+158, 
(2**17)*0+(2**8)* 48+ 71, (2**17)*0+(2**8)* 93+  3, (2**17)*1+(2**8)*119+106, 
(2**17)*0+(2**8)*  3+148, (2**17)*0+(2**8)* 53+179, (2**17)*1+(2**8)* 84+180, 
(2**17)*0+(2**8)*  5+150, (2**17)*0+(2**8)* 75+ 29, (2**17)*1+(2**8)* 75+ 70, 
(2**17)*0+(2**8)* 18+ 63, (2**17)*0+(2**8)* 40+177, (2**17)*1+(2**8)* 52+105, 
(2**17)*0+(2**8)*  8+ 14, (2**17)*0+(2**8)* 25+ 58, (2**17)*1+(2**8)* 68+127, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*0+(2**8)* 66+168, (2**17)*1+(2**8)* 69+115, 
(2**17)*0+(2**8)* 11+101, (2**17)*0+(2**8)* 14+126, (2**17)*1+(2**8)* 14+127, 
(2**17)*0+(2**8)* 10+ 63, (2**17)*0+(2**8)* 18+ 24, (2**17)*1+(2**8)* 72+ 87, 
(2**17)*0+(2**8)* 16+  7, (2**17)*0+(2**8)* 53+ 36, (2**17)*1+(2**8)* 62+ 43, 
(2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)* 18+ 44, (2**17)*1+(2**8)* 59+ 17, 
(2**17)*0+(2**8)*  4+ 50, (2**17)*0+(2**8)* 14+156, (2**17)*1+(2**8)* 72+ 12, 
(2**17)*0+(2**8)* 30+166, (2**17)*0+(2**8)* 48+ 41, (2**17)*1+(2**8)* 78+ 91, 
(2**17)*0+(2**8)*  5+ 68, (2**17)*0+(2**8)* 71+  6, (2**17)*1+(2**8)*104+ 68, 
(2**17)*0+(2**8)* 10+ 56, (2**17)*0+(2**8)* 75+115, (2**17)*1+(2**8)* 99+ 10, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*0+(2**8)* 17+ 28, (2**17)*1+(2**8)*110+ 62, 
(2**17)*0+(2**8)* 12+172, (2**17)*0+(2**8)* 18+ 84, (2**17)*1+(2**8)* 58+ 18, 
(2**17)*0+(2**8)*  7+139, (2**17)*0+(2**8)* 62+ 73, (2**17)*1+(2**8)*114+143, 
(2**17)*0+(2**8)* 12+ 33, (2**17)*0+(2**8)* 76+ 44, (2**17)*1+(2**8)* 78+ 51, 
(2**17)*0+(2**8)* 16+122, (2**17)*0+(2**8)* 60+107, (2**17)*1+(2**8)* 73+159, 
(2**17)*0+(2**8)*  2+143, (2**17)*0+(2**8)* 15+ 30, (2**17)*1+(2**8)* 87+ 26, 
(2**17)*0+(2**8)*  4+155, (2**17)*0+(2**8)* 19+106, (2**17)*1+(2**8)* 60+134, 
(2**17)*0+(2**8)* 29+ 42, (2**17)*0+(2**8)* 37+121, (2**17)*1+(2**8)* 50+ 67, 
(2**17)*0+(2**8)* 68+141, (2**17)*0+(2**8)* 71+ 68, (2**17)*1+(2**8)* 72+ 22, 
(2**17)*0+(2**8)*  3+150, (2**17)*0+(2**8)* 61+158, (2**17)*1+(2**8)*103+164, 
(2**17)*0+(2**8)* 11+131, (2**17)*0+(2**8)* 63+ 23, (2**17)*1+(2**8)* 66+ 86, 
(2**17)*0+(2**8)* 17+108, (2**17)*0+(2**8)* 70+ 16, (2**17)*1+(2**8)*110+ 78, 
(2**17)*0+(2**8)* 36+ 12, (2**17)*0+(2**8)* 80+104, (2**17)*1+(2**8)* 85+ 21, 
(2**17)*0+(2**8)*  8+ 21, (2**17)*0+(2**8)* 15+179, (2**17)*1+(2**8)* 75+167, 
(2**17)*0+(2**8)* 28+142, (2**17)*0+(2**8)* 67+ 39, (2**17)*1+(2**8)* 75+ 65, 
(2**17)*0+(2**8)* 17+ 29, (2**17)*0+(2**8)* 53+103, (2**17)*1+(2**8)* 62+107, 
(2**17)*0+(2**8)*  5+145, (2**17)*0+(2**8)* 64+ 30, (2**17)*1+(2**8)* 70+160, 
(2**17)*0+(2**8)*  2+ 69, (2**17)*0+(2**8)* 39+ 56, (2**17)*1+(2**8)* 51+137, 
(2**17)*0+(2**8)* 23+114, (2**17)*0+(2**8)* 29+ 61, (2**17)*1+(2**8)* 70+ 18, 
(2**17)*0+(2**8)*  5+ 46, (2**17)*0+(2**8)* 11+172, (2**17)*1+(2**8)* 15+143, 
(2**17)*0+(2**8)*  4+ 49, (2**17)*0+(2**8)* 10+ 70, (2**17)*1+(2**8)* 79+122, 
(2**17)*0+(2**8)* 56+ 60, (2**17)*0+(2**8)* 68+101, (2**17)*1+(2**8)* 71+ 62, 
(2**17)*0+(2**8)* 10+109, (2**17)*0+(2**8)* 75+163, (2**17)*1+(2**8)* 84+172, 
(2**17)*0+(2**8)*  4+170, (2**17)*0+(2**8)* 71+110, (2**17)*1+(2**8)* 74+163, 
(2**17)*0+(2**8)* 32+121, (2**17)*0+(2**8)* 77+  2, (2**17)*1+(2**8)* 78+ 35, 
(2**17)*0+(2**8)*  4+ 41, (2**17)*0+(2**8)* 86+146, (2**17)*1+(2**8)* 93+140, 
(2**17)*0+(2**8)* 14+ 15, (2**17)*0+(2**8)* 18+ 55, (2**17)*1+(2**8)* 63+ 58, 
(2**17)*0+(2**8)* 61+ 61, (2**17)*0+(2**8)* 66+167, (2**17)*1+(2**8)* 71+ 35, 
(2**17)*0+(2**8)* 17+ 90, (2**17)*0+(2**8)* 48+ 83, (2**17)*1+(2**8)* 63+122, 
(2**17)*0+(2**8)* 65+165, (2**17)*0+(2**8)* 67+122, (2**17)*1+(2**8)* 98+102, 
(2**17)*0+(2**8)* 37+ 22, (2**17)*0+(2**8)* 38+119, (2**17)*1+(2**8)* 56+ 92, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*0+(2**8)* 26+ 14, (2**17)*1+(2**8)* 62+ 83, 
(2**17)*0+(2**8)* 45+ 90, (2**17)*0+(2**8)* 60+156, (2**17)*1+(2**8)* 79+ 68, 
(2**17)*0+(2**8)*  4+ 72, (2**17)*0+(2**8)* 14+ 60, (2**17)*1+(2**8)* 87+120, 
(2**17)*0+(2**8)*  1+129, (2**17)*0+(2**8)*111+ 51, (2**17)*1+(2**8)*117+113, 
(2**17)*0+(2**8)* 24+ 25, (2**17)*0+(2**8)* 91+  7, (2**17)*1+(2**8)* 98+ 40, 
(2**17)*0+(2**8)* 11+119, (2**17)*0+(2**8)* 13+ 22, (2**17)*1+(2**8)* 13+ 77, 
(2**17)*0+(2**8)* 18+143, (2**17)*0+(2**8)* 35+159, (2**17)*1+(2**8)*115+134, 
(2**17)*0+(2**8)* 17+100, (2**17)*0+(2**8)* 66+ 80, (2**17)*1+(2**8)*109+147, 
(2**17)*0+(2**8)*  9+ 96, (2**17)*0+(2**8)*  9+ 12, (2**17)*1+(2**8)* 79+ 31, 
(2**17)*0+(2**8)* 12+ 65, (2**17)*0+(2**8)* 72+ 27, (2**17)*1+(2**8)* 79+109, 
(2**17)*0+(2**8)* 19+ 29, (2**17)*0+(2**8)* 79+173, (2**17)*1+(2**8)*109+112, 
(2**17)*0+(2**8)* 62+ 52, (2**17)*0+(2**8)* 63+ 84, (2**17)*1+(2**8)* 69+118, 
(2**17)*0+(2**8)* 14+ 83, (2**17)*0+(2**8)* 41+178, (2**17)*1+(2**8)* 88+176, 
(2**17)*0+(2**8)*  7+ 13, (2**17)*0+(2**8)* 41+169, (2**17)*1+(2**8)* 69+127, 
(2**17)*0+(2**8)*  0+  4, (2**17)*0+(2**8)* 14+ 84, (2**17)*1+(2**8)* 36+ 42, 
(2**17)*0+(2**8)* 61+ 64, (2**17)*0+(2**8)* 86+ 13, (2**17)*1+(2**8)* 90+ 95, 
(2**17)*0+(2**8)* 25+169, (2**17)*0+(2**8)* 70+ 64, (2**17)*1+(2**8)* 76+134, 
(2**17)*0+(2**8)* 65+148, (2**17)*0+(2**8)* 68+ 26, (2**17)*1+(2**8)* 91+ 61, 
(2**17)*0+(2**8)*  4+ 91, (2**17)*0+(2**8)*  6+ 56, (2**17)*1+(2**8)* 73+153, 
(2**17)*0+(2**8)* 13+  5, (2**17)*0+(2**8)* 39+167, (2**17)*1+(2**8)*107+  3, 
(2**17)*0+(2**8)*  9+  4, (2**17)*0+(2**8)* 66+ 59, (2**17)*1+(2**8)*102+134, 
(2**17)*0+(2**8)*  8+ 40, (2**17)*0+(2**8)* 13+ 98, (2**17)*1+(2**8)* 93+ 40, 
(2**17)*0+(2**8)*  3+ 82, (2**17)*0+(2**8)*  3+ 62, (2**17)*1+(2**8)*  6+156, 
(2**17)*0+(2**8)* 32+154, (2**17)*0+(2**8)* 45+ 28, (2**17)*1+(2**8)* 88+171, 
(2**17)*0+(2**8)*  6+ 65, (2**17)*0+(2**8)* 55+122, (2**17)*1+(2**8)*102+159, 
(2**17)*0+(2**8)*  0+145, (2**17)*0+(2**8)* 16+147, (2**17)*1+(2**8)*100+ 90, 
(2**17)*0+(2**8)* 61+ 78, (2**17)*0+(2**8)* 68+ 48, (2**17)*1+(2**8)*116+ 11, 
(2**17)*0+(2**8)*  1+ 62, (2**17)*0+(2**8)* 62+  7, (2**17)*1+(2**8)* 69+ 47, 
(2**17)*0+(2**8)* 19+ 76, (2**17)*0+(2**8)* 52+162, (2**17)*1+(2**8)* 72+ 58, 
(2**17)*0+(2**8)* 43+174, (2**17)*0+(2**8)* 69+ 62, (2**17)*1+(2**8)* 72+ 52, 
(2**17)*0+(2**8)* 20+166, (2**17)*0+(2**8)*107+147, (2**17)*1+(2**8)*118+109, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*0+(2**8)* 17+176, (2**17)*1+(2**8)* 73+101, 
(2**17)*0+(2**8)*  7+119, (2**17)*0+(2**8)* 75+ 54, (2**17)*1+(2**8)*109+ 35, 
(2**17)*0+(2**8)* 17+ 49, (2**17)*0+(2**8)* 74+166, (2**17)*1+(2**8)* 94+ 54, 
(2**17)*0+(2**8)*  4+121, (2**17)*0+(2**8)* 19+142, (2**17)*1+(2**8)* 79+145, 
(2**17)*0+(2**8)* 16+166, (2**17)*0+(2**8)* 21+162, (2**17)*1+(2**8)* 91+ 65, 
(2**17)*0+(2**8)* 21+ 59, (2**17)*0+(2**8)* 40+ 28, (2**17)*1+(2**8)* 73+174, 
(2**17)*0+(2**8)* 72+ 99, (2**17)*0+(2**8)* 90+174, (2**17)*1+(2**8)*111+ 21, 
(2**17)*0+(2**8)*  1+ 48, (2**17)*0+(2**8)*  5+ 36, (2**17)*1+(2**8)*  7+  5, 
(2**17)*0+(2**8)*  3+ 88, (2**17)*0+(2**8)* 42+131, (2**17)*1+(2**8)* 63+ 34, 
(2**17)*0+(2**8)*  1+ 28, (2**17)*0+(2**8)*  7+ 25, (2**17)*1+(2**8)*  8+ 81, 
(2**17)*0+(2**8)*  2+148, (2**17)*0+(2**8)* 74+123, (2**17)*1+(2**8)* 96+152, 
(2**17)*0+(2**8)* 44+156, (2**17)*0+(2**8)* 60+ 23, (2**17)*1+(2**8)* 60+ 88, 
(2**17)*0+(2**8)* 95+114, (2**17)*0+(2**8)*106+ 92, (2**17)*1+(2**8)*114+118, 
(2**17)*0+(2**8)*  6+ 71, (2**17)*0+(2**8)* 16+121, (2**17)*1+(2**8)* 87+142, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*0+(2**8)* 46+104, (2**17)*1+(2**8)* 72+166, 
(2**17)*0+(2**8)* 10+177, (2**17)*0+(2**8)* 23+172, (2**17)*1+(2**8)* 73+ 10, 
(2**17)*0+(2**8)*  4+100, (2**17)*0+(2**8)* 77+ 43, (2**17)*1+(2**8)* 78+  8, 
(2**17)*0+(2**8)*  5+ 51, (2**17)*0+(2**8)*  5+ 94, (2**17)*1+(2**8)* 15+131, 
(2**17)*0+(2**8)*  9+ 50, (2**17)*0+(2**8)* 47+ 33, (2**17)*1+(2**8)* 78+ 64, 
(2**17)*0+(2**8)* 21+ 72, (2**17)*0+(2**8)* 22+ 66, (2**17)*1+(2**8)* 94+165, 
(2**17)*0+(2**8)*  9+144, (2**17)*0+(2**8)* 23+113, (2**17)*1+(2**8)* 76+ 27, 
(2**17)*0+(2**8)*  2+ 48, (2**17)*0+(2**8)* 19+ 88, (2**17)*1+(2**8)* 45+131, 
(2**17)*0+(2**8)*  9+ 31, (2**17)*0+(2**8)* 68+156, (2**17)*1+(2**8)* 76+ 54, 
(2**17)*0+(2**8)* 14+ 75, (2**17)*0+(2**8)* 16+155, (2**17)*1+(2**8)* 54+ 20, 
(2**17)*0+(2**8)* 60+ 67, (2**17)*0+(2**8)* 70+ 72, (2**17)*1+(2**8)* 71+ 31, 
(2**17)*0+(2**8)*  0+ 68, (2**17)*0+(2**8)* 22+161, (2**17)*1+(2**8)* 62+112, 
(2**17)*0+(2**8)* 44+ 59, (2**17)*0+(2**8)* 67+164, (2**17)*1+(2**8)* 71+ 46, 
(2**17)*0+(2**8)* 77+  3, (2**17)*0+(2**8)*112+  5, (2**17)*1+(2**8)*117+ 33, 
(2**17)*0+(2**8)* 13+118, (2**17)*0+(2**8)* 35+122, (2**17)*1+(2**8)* 94+ 88, 
(2**17)*0+(2**8)*  7+130, (2**17)*0+(2**8)* 68+103, (2**17)*1+(2**8)*118+ 44, 
(2**17)*0+(2**8)* 22+118, (2**17)*0+(2**8)* 46+105, (2**17)*1+(2**8)* 70+163, 
(2**17)*0+(2**8)* 10+ 48, (2**17)*0+(2**8)* 14+ 31, (2**17)*1+(2**8)* 92+166, 
(2**17)*0+(2**8)*  5+169, (2**17)*0+(2**8)* 11+ 97, (2**17)*1+(2**8)* 76+119, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*0+(2**8)*  7+ 80, (2**17)*1+(2**8)* 12+138, 
(2**17)*0+(2**8)* 17+ 36, (2**17)*0+(2**8)* 63+ 33, (2**17)*1+(2**8)* 89+ 74, 
(2**17)*0+(2**8)* 43+ 77, (2**17)*0+(2**8)* 69+ 96, (2**17)*1+(2**8)* 97+ 80, 
(2**17)*0+(2**8)*  6+ 18, (2**17)*0+(2**8)* 75+ 79, (2**17)*1+(2**8)* 78+119, 
(2**17)*0+(2**8)* 60+  2, (2**17)*0+(2**8)* 65+ 83, (2**17)*1+(2**8)* 68+127, 
(2**17)*0+(2**8)*  2+ 53, (2**17)*0+(2**8)* 67+149, (2**17)*1+(2**8)*115+ 17, 
(2**17)*0+(2**8)*  4+106, (2**17)*0+(2**8)* 57+161, (2**17)*1+(2**8)* 77+ 48, 
(2**17)*0+(2**8)* 13+ 93, (2**17)*0+(2**8)* 20+117, (2**17)*1+(2**8)*101+107, 
(2**17)*0+(2**8)* 16+ 72, (2**17)*0+(2**8)* 61+137, (2**17)*1+(2**8)* 66+169, 
(2**17)*0+(2**8)*  4+149, (2**17)*0+(2**8)* 13+143, (2**17)*1+(2**8)* 59+165, 
(2**17)*0+(2**8)* 19+157, (2**17)*0+(2**8)* 65+121, (2**17)*1+(2**8)* 66+  7, 
(2**17)*0+(2**8)* 33+  2, (2**17)*0+(2**8)* 59+105, (2**17)*1+(2**8)*108+ 71, 
(2**17)*0+(2**8)* 24+179, (2**17)*0+(2**8)* 63+148, (2**17)*1+(2**8)*113+179, 
(2**17)*0+(2**8)* 15+ 28, (2**17)*0+(2**8)* 15+ 69, (2**17)*1+(2**8)* 65+150, 
(2**17)*0+(2**8)* 78+ 63, (2**17)*0+(2**8)*100+177, (2**17)*1+(2**8)*112+105, 
(2**17)*0+(2**8)*  8+126, (2**17)*0+(2**8)* 68+ 14, (2**17)*1+(2**8)* 85+ 58, 
(2**17)*0+(2**8)*  6+167, (2**17)*0+(2**8)*  9+114, (2**17)*1+(2**8)* 60+ 77, 
(2**17)*0+(2**8)* 71+101, (2**17)*0+(2**8)* 74+126, (2**17)*1+(2**8)* 74+127, 
(2**17)*0+(2**8)* 12+ 86, (2**17)*0+(2**8)* 70+ 63, (2**17)*1+(2**8)* 78+ 24, 
(2**17)*0+(2**8)*  2+ 42, (2**17)*0+(2**8)* 76+  7, (2**17)*1+(2**8)*113+ 36, 
(2**17)*0+(2**8)* 67+ 51, (2**17)*0+(2**8)* 78+ 44, (2**17)*1+(2**8)*119+ 17, 
(2**17)*0+(2**8)* 12+ 11, (2**17)*0+(2**8)* 64+ 50, (2**17)*1+(2**8)* 74+156, 
(2**17)*0+(2**8)* 18+ 90, (2**17)*0+(2**8)* 90+166, (2**17)*1+(2**8)*108+ 41, 
(2**17)*0+(2**8)* 11+  5, (2**17)*0+(2**8)* 44+ 67, (2**17)*1+(2**8)* 65+ 68, 
(2**17)*0+(2**8)* 15+114, (2**17)*0+(2**8)* 39+  9, (2**17)*1+(2**8)* 70+ 56, 
(2**17)*0+(2**8)* 50+ 61, (2**17)*0+(2**8)* 60+ 87, (2**17)*1+(2**8)* 77+ 28, 
(2**17)*0+(2**8)* 72+172, (2**17)*0+(2**8)* 78+ 84, (2**17)*1+(2**8)*118+ 18, 
(2**17)*0+(2**8)*  2+ 72, (2**17)*0+(2**8)* 54+142, (2**17)*1+(2**8)* 67+139, 
(2**17)*0+(2**8)* 16+ 43, (2**17)*0+(2**8)* 18+ 50, (2**17)*1+(2**8)* 72+ 33, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)* 13+158, (2**17)*1+(2**8)* 76+122, 
(2**17)*0+(2**8)* 27+ 25, (2**17)*0+(2**8)* 62+143, (2**17)*1+(2**8)* 75+ 30, 
(2**17)*0+(2**8)*  0+133, (2**17)*0+(2**8)* 64+155, (2**17)*1+(2**8)* 79+106, 
(2**17)*0+(2**8)* 89+ 42, (2**17)*0+(2**8)* 97+121, (2**17)*1+(2**8)*110+ 67, 
(2**17)*0+(2**8)*  8+140, (2**17)*0+(2**8)* 11+ 67, (2**17)*1+(2**8)* 12+ 21, 
(2**17)*0+(2**8)*  1+157, (2**17)*0+(2**8)* 43+163, (2**17)*1+(2**8)* 63+150, 
(2**17)*0+(2**8)*  3+ 22, (2**17)*0+(2**8)*  6+ 85, (2**17)*1+(2**8)* 71+131, 
(2**17)*0+(2**8)* 10+ 15, (2**17)*0+(2**8)* 50+ 77, (2**17)*1+(2**8)* 77+108, 
(2**17)*0+(2**8)* 20+103, (2**17)*0+(2**8)* 25+ 20, (2**17)*1+(2**8)* 96+ 12, 
(2**17)*0+(2**8)* 15+166, (2**17)*0+(2**8)* 68+ 21, (2**17)*1+(2**8)* 75+179, 
(2**17)*0+(2**8)*  7+ 38, (2**17)*0+(2**8)* 15+ 64, (2**17)*1+(2**8)* 88+142, 
(2**17)*0+(2**8)*  2+106, (2**17)*0+(2**8)* 77+ 29, (2**17)*1+(2**8)*113+103, 
(2**17)*0+(2**8)*  4+ 29, (2**17)*0+(2**8)* 10+159, (2**17)*1+(2**8)* 65+145, 
(2**17)*0+(2**8)* 62+ 69, (2**17)*0+(2**8)* 99+ 56, (2**17)*1+(2**8)*111+137, 
(2**17)*0+(2**8)* 10+ 17, (2**17)*0+(2**8)* 83+114, (2**17)*1+(2**8)* 89+ 61, 
(2**17)*0+(2**8)* 65+ 46, (2**17)*0+(2**8)* 71+172, (2**17)*1+(2**8)* 75+143, 
(2**17)*0+(2**8)* 19+121, (2**17)*0+(2**8)* 64+ 49, (2**17)*1+(2**8)* 70+ 70, 
(2**17)*0+(2**8)*  8+100, (2**17)*0+(2**8)* 11+ 61, (2**17)*1+(2**8)*116+ 60, 
(2**17)*0+(2**8)* 15+162, (2**17)*0+(2**8)* 24+171, (2**17)*1+(2**8)* 70+109, 
(2**17)*0+(2**8)* 11+109, (2**17)*0+(2**8)* 14+162, (2**17)*1+(2**8)* 64+170, 
(2**17)*0+(2**8)* 17+  1, (2**17)*0+(2**8)* 18+ 34, (2**17)*1+(2**8)* 92+121, 
(2**17)*0+(2**8)* 26+145, (2**17)*0+(2**8)* 33+139, (2**17)*1+(2**8)* 64+ 41, 
(2**17)*0+(2**8)*  3+ 57, (2**17)*0+(2**8)* 74+ 15, (2**17)*1+(2**8)* 78+ 55, 
(2**17)*0+(2**8)*  1+ 60, (2**17)*0+(2**8)*  6+166, (2**17)*1+(2**8)* 11+ 34, 
(2**17)*0+(2**8)*  3+121, (2**17)*0+(2**8)* 77+ 90, (2**17)*1+(2**8)*108+ 83, 
(2**17)*0+(2**8)*  5+164, (2**17)*0+(2**8)*  7+121, (2**17)*1+(2**8)* 38+101, 
(2**17)*0+(2**8)* 97+ 22, (2**17)*0+(2**8)* 98+119, (2**17)*1+(2**8)*116+ 92, 
(2**17)*0+(2**8)*  2+ 82, (2**17)*0+(2**8)* 61+ 92, (2**17)*1+(2**8)* 86+ 14, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)* 19+ 67, (2**17)*1+(2**8)*105+ 90, 
(2**17)*0+(2**8)* 27+119, (2**17)*0+(2**8)* 64+ 72, (2**17)*1+(2**8)* 74+ 60, 
(2**17)*0+(2**8)* 51+ 50, (2**17)*0+(2**8)* 57+112, (2**17)*1+(2**8)* 61+129, 
(2**17)*0+(2**8)* 31+  6, (2**17)*0+(2**8)* 38+ 39, (2**17)*1+(2**8)* 84+ 25, 
(2**17)*0+(2**8)* 71+119, (2**17)*0+(2**8)* 73+ 22, (2**17)*1+(2**8)* 73+ 77, 
(2**17)*0+(2**8)* 55+133, (2**17)*0+(2**8)* 78+143, (2**17)*1+(2**8)* 95+159, 
(2**17)*0+(2**8)*  6+ 79, (2**17)*0+(2**8)* 49+146, (2**17)*1+(2**8)* 77+100, 
(2**17)*0+(2**8)* 19+ 30, (2**17)*0+(2**8)* 69+ 96, (2**17)*1+(2**8)* 69+ 12, 
(2**17)*0+(2**8)* 12+ 26, (2**17)*0+(2**8)* 19+108, (2**17)*1+(2**8)* 72+ 65, 
(2**17)*0+(2**8)* 19+172, (2**17)*0+(2**8)* 49+111, (2**17)*1+(2**8)* 79+ 29, 
(2**17)*0+(2**8)*  2+ 51, (2**17)*0+(2**8)*  3+ 83, (2**17)*1+(2**8)*  9+117, 
(2**17)*0+(2**8)* 28+175, (2**17)*0+(2**8)* 74+ 83, (2**17)*1+(2**8)*101+178, 
(2**17)*0+(2**8)*  9+126, (2**17)*0+(2**8)* 67+ 13, (2**17)*1+(2**8)*101+169, 
(2**17)*0+(2**8)* 60+  4, (2**17)*0+(2**8)* 74+ 84, (2**17)*1+(2**8)* 96+ 42, 
(2**17)*0+(2**8)*  1+ 63, (2**17)*0+(2**8)* 26+ 12, (2**17)*1+(2**8)* 30+ 94, 
(2**17)*0+(2**8)* 10+ 63, (2**17)*0+(2**8)* 16+133, (2**17)*1+(2**8)* 85+169, 
(2**17)*0+(2**8)*  5+147, (2**17)*0+(2**8)*  8+ 25, (2**17)*1+(2**8)* 31+ 60, 
(2**17)*0+(2**8)* 13+152, (2**17)*0+(2**8)* 64+ 91, (2**17)*1+(2**8)* 66+ 56, 
(2**17)*0+(2**8)* 47+  2, (2**17)*0+(2**8)* 73+  5, (2**17)*1+(2**8)* 99+167, 
(2**17)*0+(2**8)*  6+ 58, (2**17)*0+(2**8)* 42+133, (2**17)*1+(2**8)* 69+  4, 
(2**17)*0+(2**8)* 33+ 39, (2**17)*0+(2**8)* 68+ 40, (2**17)*1+(2**8)* 73+ 98, 
(2**17)*0+(2**8)* 63+ 82, (2**17)*0+(2**8)* 63+ 62, (2**17)*1+(2**8)* 66+156, 
(2**17)*0+(2**8)* 28+170, (2**17)*0+(2**8)* 92+154, (2**17)*1+(2**8)*105+ 28, 
(2**17)*0+(2**8)* 42+158, (2**17)*0+(2**8)* 66+ 65, (2**17)*1+(2**8)*115+122, 
(2**17)*0+(2**8)* 40+ 89, (2**17)*0+(2**8)* 60+145, (2**17)*1+(2**8)* 76+147, 
(2**17)*0+(2**8)*  1+ 77, (2**17)*0+(2**8)*  8+ 47, (2**17)*1+(2**8)* 56+ 10, 
(2**17)*0+(2**8)*  2+  6, (2**17)*0+(2**8)*  9+ 46, (2**17)*1+(2**8)* 61+ 62, 
(2**17)*0+(2**8)* 12+ 57, (2**17)*0+(2**8)* 79+ 76, (2**17)*1+(2**8)*112+162, 
(2**17)*0+(2**8)*  9+ 61, (2**17)*0+(2**8)* 12+ 51, (2**17)*1+(2**8)*103+174, 
(2**17)*0+(2**8)* 47+146, (2**17)*0+(2**8)* 58+108, (2**17)*1+(2**8)* 80+166, 
(2**17)*0+(2**8)* 13+100, (2**17)*0+(2**8)* 63+ 83, (2**17)*1+(2**8)* 77+176, 
(2**17)*0+(2**8)* 15+ 53, (2**17)*0+(2**8)* 49+ 34, (2**17)*1+(2**8)* 67+119, 
(2**17)*0+(2**8)* 14+165, (2**17)*0+(2**8)* 34+ 53, (2**17)*1+(2**8)* 77+ 49, 
(2**17)*0+(2**8)* 19+144, (2**17)*0+(2**8)* 64+121, (2**17)*1+(2**8)* 79+142, 
(2**17)*0+(2**8)* 31+ 64, (2**17)*0+(2**8)* 76+166, (2**17)*1+(2**8)* 81+162, 
(2**17)*0+(2**8)* 13+173, (2**17)*0+(2**8)* 81+ 59, (2**17)*1+(2**8)*100+ 28, 
(2**17)*0+(2**8)* 12+ 98, (2**17)*0+(2**8)* 30+173, (2**17)*1+(2**8)* 51+ 20, 
(2**17)*0+(2**8)* 61+ 48, (2**17)*0+(2**8)* 65+ 36, (2**17)*1+(2**8)* 67+  5, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*0+(2**8)* 63+ 88, (2**17)*1+(2**8)*102+131, 
(2**17)*0+(2**8)* 61+ 28, (2**17)*0+(2**8)* 67+ 25, (2**17)*1+(2**8)* 68+ 81, 
(2**17)*0+(2**8)* 14+122, (2**17)*0+(2**8)* 36+151, (2**17)*1+(2**8)* 62+148, 


(2**17)*0+(2**8)*  0+ 23, (2**17)*0+(2**8)*  0+ 88, (2**17)*0+(2**8)* 71+142, (2**17)*1+(2**8)*104+132, 
(2**17)*0+(2**8)* 19+ 64, (2**17)*0+(2**8)* 45+ 33, (2**17)*0+(2**8)* 89+122, (2**17)*1+(2**8)* 95+ 87, 
(2**17)*0+(2**8)*  6+156, (2**17)*0+(2**8)* 28+107, (2**17)*0+(2**8)* 83+178, (2**17)*1+(2**8)*112+ 69, 
(2**17)*0+(2**8)* 49+149, (2**17)*0+(2**8)* 73+ 64, (2**17)*0+(2**8)* 84+156, (2**17)*1+(2**8)* 95+107, 
(2**17)*0+(2**8)* 13+166, (2**17)*0+(2**8)* 77+ 95, (2**17)*0+(2**8)* 88+132, (2**17)*1+(2**8)*143+ 69, 
(2**17)*0+(2**8)* 14+ 10, (2**17)*0+(2**8)* 66+157, (2**17)*0+(2**8)* 76+101, (2**17)*1+(2**8)* 77+ 52, 
(2**17)*0+(2**8)* 17+ 27, (2**17)*0+(2**8)* 44+ 75, (2**17)*0+(2**8)* 82+115, (2**17)*1+(2**8)* 89+125, 
(2**17)*0+(2**8)*  9+156, (2**17)*0+(2**8)* 24+ 80, (2**17)*0+(2**8)*104+ 31, (2**17)*1+(2**8)*133+159, 
(2**17)*0+(2**8)* 46+ 44, (2**17)*0+(2**8)* 80+112, (2**17)*0+(2**8)* 84+ 68, (2**17)*1+(2**8)* 92+ 89, 
(2**17)*0+(2**8)* 10+  4, (2**17)*0+(2**8)* 43+140, (2**17)*0+(2**8)* 74+ 49, (2**17)*1+(2**8)* 91+110, 
(2**17)*0+(2**8)* 11+ 72, (2**17)*0+(2**8)* 18+113, (2**17)*0+(2**8)* 21+115, (2**17)*1+(2**8)*139+ 50, 
(2**17)*0+(2**8)* 12+ 31, (2**17)*0+(2**8)* 15+ 83, (2**17)*0+(2**8)* 17+ 54, (2**17)*1+(2**8)* 42+ 80, 
(2**17)*0+(2**8)*  0+ 67, (2**17)*0+(2**8)*  2+112, (2**17)*0+(2**8)* 21+ 19, (2**17)*1+(2**8)*118+102, 
(2**17)*0+(2**8)*  7+164, (2**17)*0+(2**8)* 72+ 69, (2**17)*0+(2**8)* 80+155, (2**17)*1+(2**8)*132+103, 
(2**17)*0+(2**8)* 86+119, (2**17)*0+(2**8)* 98+145, (2**17)*0+(2**8)* 99+155, (2**17)*1+(2**8)*119+109, 
(2**17)*0+(2**8)* 22+132, (2**17)*0+(2**8)* 23+177, (2**17)*0+(2**8)* 57+ 61, (2**17)*1+(2**8)* 86+102, 
(2**17)*0+(2**8)* 17+119, (2**17)*0+(2**8)* 21+ 93, (2**17)*0+(2**8)* 87+123, (2**17)*1+(2**8)*131+ 49, 
(2**17)*0+(2**8)*  8+162, (2**17)*0+(2**8)* 23+114, (2**17)*0+(2**8)* 76+ 60, (2**17)*1+(2**8)*131+  6, 
(2**17)*0+(2**8)*  9+103, (2**17)*0+(2**8)* 21+ 56, (2**17)*0+(2**8)* 63+ 98, (2**17)*1+(2**8)* 79+ 81, 
(2**17)*0+(2**8)*  8+107, (2**17)*0+(2**8)* 11+163, (2**17)*0+(2**8)* 68+ 61, (2**17)*1+(2**8)* 78+168, 
(2**17)*0+(2**8)*  5+ 83, (2**17)*0+(2**8)* 59+  7, (2**17)*0+(2**8)* 73+158, (2**17)*1+(2**8)* 85+139, 
(2**17)*0+(2**8)*  7+149, (2**17)*0+(2**8)* 86+144, (2**17)*0+(2**8)* 94+  7, (2**17)*1+(2**8)*120+ 87, 
(2**17)*0+(2**8)* 16+ 26, (2**17)*0+(2**8)* 56+ 35, (2**17)*0+(2**8)* 74+ 54, (2**17)*1+(2**8)* 84+ 98, 
(2**17)*0+(2**8)*  0+  2, (2**17)*0+(2**8)*  9+127, (2**17)*0+(2**8)* 65+ 92, (2**17)*1+(2**8)* 82+ 47, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*0+(2**8)*  4+ 37, (2**17)*0+(2**8)*  5+121, (2**17)*1+(2**8)* 49+127, 
(2**17)*0+(2**8)* 16+ 79, (2**17)*0+(2**8)* 19+ 63, (2**17)*0+(2**8)* 24+ 88, (2**17)*1+(2**8)* 56+ 49, 
(2**17)*0+(2**8)* 76+107, (2**17)*0+(2**8)* 80+ 71, (2**17)*0+(2**8)* 91+ 52, (2**17)*1+(2**8)*125+133, 
(2**17)*0+(2**8)*  1+137, (2**17)*0+(2**8)* 39+117, (2**17)*0+(2**8)* 88+ 29, (2**17)*1+(2**8)* 94+143, 
(2**17)*0+(2**8)*  8+ 80, (2**17)*0+(2**8)* 78+167, (2**17)*0+(2**8)*106+ 38, (2**17)*1+(2**8)*122+140, 
(2**17)*0+(2**8)* 23+ 12, (2**17)*0+(2**8)* 73+ 77, (2**17)*0+(2**8)* 76+150, (2**17)*1+(2**8)*136+165, 
(2**17)*0+(2**8)*  3+ 88, (2**17)*0+(2**8)* 78+ 86, (2**17)*0+(2**8)* 90+165, (2**17)*1+(2**8)*123+130, 
(2**17)*0+(2**8)* 11+ 90, (2**17)*0+(2**8)* 27+177, (2**17)*0+(2**8)* 53+ 91, (2**17)*1+(2**8)* 78+ 72, 
(2**17)*0+(2**8)* 38+ 67, (2**17)*0+(2**8)* 81+ 17, (2**17)*0+(2**8)* 87+ 32, (2**17)*1+(2**8)* 90+ 52, 
(2**17)*0+(2**8)* 69+144, (2**17)*0+(2**8)* 81+127, (2**17)*0+(2**8)* 89+ 73, (2**17)*1+(2**8)*103+105, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*0+(2**8)* 10+ 96, (2**17)*0+(2**8)* 15+156, (2**17)*1+(2**8)* 57+124, 
(2**17)*0+(2**8)*  6+ 56, (2**17)*0+(2**8)* 13+ 50, (2**17)*0+(2**8)* 67+131, (2**17)*1+(2**8)* 93+114, 
(2**17)*0+(2**8)*  9+ 14, (2**17)*0+(2**8)* 87+166, (2**17)*0+(2**8)* 89+ 44, (2**17)*1+(2**8)*120+133, 
(2**17)*0+(2**8)* 11+ 63, (2**17)*0+(2**8)* 74+ 43, (2**17)*0+(2**8)*105+136, (2**17)*1+(2**8)*137+ 54, 
(2**17)*0+(2**8)* 12+101, (2**17)*0+(2**8)* 13+172, (2**17)*0+(2**8)* 80+ 78, (2**17)*1+(2**8)*134+ 62, 
(2**17)*0+(2**8)*  4+ 50, (2**17)*0+(2**8)* 37+ 39, (2**17)*0+(2**8)* 83+ 72, (2**17)*1+(2**8)* 85+ 87, 
(2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)* 88+ 70, (2**17)*0+(2**8)* 94+ 61, (2**17)*1+(2**8)*122+147, 
(2**17)*0+(2**8)*  4+155, (2**17)*0+(2**8)*  5+ 68, (2**17)*0+(2**8)* 91+ 91, (2**17)*1+(2**8)*122+131, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*0+(2**8)* 13+131, (2**17)*0+(2**8)* 90+ 53, (2**17)*1+(2**8)*130+170, 
(2**17)*0+(2**8)* 11+ 56, (2**17)*0+(2**8)* 25+147, (2**17)*0+(2**8)* 68+101, (2**17)*1+(2**8)* 90+128, 
(2**17)*0+(2**8)*  7+139, (2**17)*0+(2**8)* 16+179, (2**17)*0+(2**8)* 69+ 20, (2**17)*1+(2**8)* 87+ 81, 
(2**17)*0+(2**8)*  2+115, (2**17)*0+(2**8)* 37+120, (2**17)*0+(2**8)* 83+ 16, (2**17)*1+(2**8)* 85+ 12, 
(2**17)*0+(2**8)* 23+159, (2**17)*0+(2**8)* 72+107, (2**17)*0+(2**8)*104+  5, (2**17)*1+(2**8)*130+ 74, 
(2**17)*0+(2**8)* 19+ 24, (2**17)*0+(2**8)* 78+ 33, (2**17)*0+(2**8)* 86+159, (2**17)*1+(2**8)*140+ 98, 
(2**17)*0+(2**8)*  2+143, (2**17)*0+(2**8)* 41+ 36, (2**17)*0+(2**8)* 72+134, (2**17)*1+(2**8)* 93+173, 
(2**17)*0+(2**8)* 75+ 34, (2**17)*0+(2**8)* 83+160, (2**17)*0+(2**8)* 92+158, (2**17)*1+(2**8)*109+ 62, 
(2**17)*0+(2**8)*  1+ 62, (2**17)*0+(2**8)* 23+ 42, (2**17)*0+(2**8)* 75+ 84, (2**17)*1+(2**8)*124+ 62, 
(2**17)*0+(2**8)* 75+101, (2**17)*0+(2**8)* 85+ 22, (2**17)*0+(2**8)*106+ 94, (2**17)*1+(2**8)*116+ 10, 
(2**17)*0+(2**8)* 12+172, (2**17)*0+(2**8)* 27+115, (2**17)*0+(2**8)* 69+ 22, (2**17)*1+(2**8)* 81+141, 
(2**17)*0+(2**8)* 17+122, (2**17)*0+(2**8)* 90+ 33, (2**17)*0+(2**8)* 94+ 65, (2**17)*1+(2**8)*134+164, 
(2**17)*0+(2**8)*  6+  7, (2**17)*0+(2**8)*  9+ 21, (2**17)*0+(2**8)* 13+ 33, (2**17)*1+(2**8)* 38+ 91, 
(2**17)*0+(2**8)*  8+104, (2**17)*0+(2**8)* 18+175, (2**17)*0+(2**8)* 19+ 84, (2**17)*1+(2**8)* 57+ 48, 
(2**17)*0+(2**8)*  8+ 24, (2**17)*0+(2**8)* 25+ 56, (2**17)*0+(2**8)* 52+ 58, (2**17)*1+(2**8)* 79+ 39, 
(2**17)*0+(2**8)* 22+166, (2**17)*0+(2**8)* 84+110, (2**17)*0+(2**8)* 88+163, (2**17)*1+(2**8)*136+ 81, 
(2**17)*0+(2**8)*  2+ 69, (2**17)*0+(2**8)* 10+145, (2**17)*0+(2**8)* 47+156, (2**17)*1+(2**8)* 74+107, 
(2**17)*0+(2**8)* 51+ 39, (2**17)*0+(2**8)* 81+101, (2**17)*0+(2**8)* 84+ 35, (2**17)*1+(2**8)*107+124, 
(2**17)*0+(2**8)*  5+145, (2**17)*0+(2**8)* 33+ 92, (2**17)*0+(2**8)* 83+ 18, (2**17)*1+(2**8)*113+  6, 
(2**17)*0+(2**8)* 11+ 70, (2**17)*0+(2**8)* 20+106, (2**17)*0+(2**8)* 86+143, (2**17)*1+(2**8)*118+180, 
(2**17)*0+(2**8)*  4+ 49, (2**17)*0+(2**8)* 40+118, (2**17)*0+(2**8)* 78+ 19, (2**17)*1+(2**8)* 95+100, 
(2**17)*0+(2**8)* 19+ 55, (2**17)*0+(2**8)* 90+160, (2**17)*0+(2**8)* 94+177, (2**17)*1+(2**8)*138+156, 
(2**17)*0+(2**8)*  4+170, (2**17)*0+(2**8)*  5+ 46, (2**17)*0+(2**8)* 91+ 35, (2**17)*1+(2**8)*117+ 91, 
(2**17)*0+(2**8)* 77+165, (2**17)*0+(2**8)* 88+167, (2**17)*0+(2**8)*101+168, (2**17)*1+(2**8)*123+ 71, 
(2**17)*0+(2**8)* 58+ 99, (2**17)*0+(2**8)* 75+ 58, (2**17)*0+(2**8)* 84+ 62, (2**17)*1+(2**8)* 88+ 65, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*0+(2**8)*  8+ 95, (2**17)*0+(2**8)*102+  1, (2**17)*1+(2**8)*108+138, 
(2**17)*0+(2**8)*  4+ 72, (2**17)*0+(2**8)* 33+ 16, (2**17)*0+(2**8)* 88+169, (2**17)*1+(2**8)*114+143, 
(2**17)*0+(2**8)* 35+168, (2**17)*0+(2**8)* 49+105, (2**17)*0+(2**8)* 79+122, (2**17)*1+(2**8)* 91+ 51, 
(2**17)*0+(2**8)*  8+  3, (2**17)*0+(2**8)* 73+ 62, (2**17)*0+(2**8)* 91+165, (2**17)*1+(2**8)*114+ 25, 
(2**17)*0+(2**8)* 11+109, (2**17)*0+(2**8)* 23+ 27, (2**17)*0+(2**8)* 72+156, (2**17)*1+(2**8)*126+ 21, 
(2**17)*0+(2**8)* 18+ 82, (2**17)*0+(2**8)* 55+ 55, (2**17)*0+(2**8)* 74+ 83, (2**17)*1+(2**8)* 93+119, 
(2**17)*0+(2**8)* 43+125, (2**17)*0+(2**8)* 73+ 78, (2**17)*0+(2**8)* 80+ 25, (2**17)*1+(2**8)* 92+122, 
(2**17)*0+(2**8)* 12+119, (2**17)*0+(2**8)* 12+ 46, (2**17)*0+(2**8)*103+ 68, (2**17)*1+(2**8)*125+ 12, 
(2**17)*0+(2**8)* 30+ 33, (2**17)*0+(2**8)* 90+ 37, (2**17)*0+(2**8)*101+ 49, (2**17)*1+(2**8)*120+ 84, 
(2**17)*0+(2**8)* 15+126, (2**17)*0+(2**8)* 24+126, (2**17)*0+(2**8)* 38+170, (2**17)*1+(2**8)* 75+115, 
(2**17)*0+(2**8)* 22+150, (2**17)*0+(2**8)* 93+ 67, (2**17)*0+(2**8)*103+177, (2**17)*1+(2**8)*142+ 26, 
(2**17)*0+(2**8)* 14+ 77, (2**17)*0+(2**8)* 70+ 22, (2**17)*0+(2**8)* 82+ 32, (2**17)*1+(2**8)* 85+ 27, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*0+(2**8)* 12+131, (2**17)*0+(2**8)* 71+ 78, (2**17)*1+(2**8)* 90+175, 
(2**17)*0+(2**8)*  7+ 13, (2**17)*0+(2**8)*  7+172, (2**17)*0+(2**8)* 74+ 52, (2**17)*1+(2**8)*133+ 24, 
(2**17)*0+(2**8)* 10+ 12, (2**17)*0+(2**8)* 19+143, (2**17)*0+(2**8)* 94+ 40, (2**17)*1+(2**8)*135+  7, 
(2**17)*0+(2**8)* 92+ 31, (2**17)*0+(2**8)* 92+109, (2**17)*0+(2**8)* 95+152, (2**17)*1+(2**8)*111+ 34, 
(2**17)*0+(2**8)*  0+  4, (2**17)*0+(2**8)* 77+148, (2**17)*0+(2**8)* 82+118, (2**17)*1+(2**8)*139+ 93, 
(2**17)*0+(2**8)*  1+ 28, (2**17)*0+(2**8)* 20+ 29, (2**17)*0+(2**8)* 92+173, (2**17)*1+(2**8)*124+ 69, 
(2**17)*0+(2**8)*  6+ 65, (2**17)*0+(2**8)* 18+100, (2**17)*0+(2**8)* 65+153, (2**17)*1+(2**8)* 82+127, 
(2**17)*0+(2**8)* 10+ 32, (2**17)*0+(2**8)* 86+153, (2**17)*0+(2**8)* 87+ 76, (2**17)*1+(2**8)*132+169, 
(2**17)*0+(2**8)* 20+ 93, (2**17)*0+(2**8)* 66+ 36, (2**17)*0+(2**8)* 89+134, (2**17)*1+(2**8)*100+176, 
(2**17)*0+(2**8)*  4+ 91, (2**17)*0+(2**8)* 26+ 56, (2**17)*0+(2**8)* 81+ 26, (2**17)*1+(2**8)*108+ 63, 
(2**17)*0+(2**8)* 23+126, (2**17)*0+(2**8)* 78+ 59, (2**17)*0+(2**8)* 82+ 51, (2**17)*1+(2**8)*127+ 39, 
(2**17)*0+(2**8)*  3+150, (2**17)*0+(2**8)*  6+169, (2**17)*0+(2**8)* 55+131, (2**17)*1+(2**8)* 87+107, 
(2**17)*0+(2**8)*  3+ 62, (2**17)*0+(2**8)* 14+ 98, (2**17)*0+(2**8)*102+164, (2**17)*1+(2**8)*108+ 35, 
(2**17)*0+(2**8)*  5+154, (2**17)*0+(2**8)*  9+ 40, (2**17)*0+(2**8)* 25+119, (2**17)*1+(2**8)*126+122, 
(2**17)*0+(2**8)*  0+145, (2**17)*0+(2**8)* 22+ 99, (2**17)*0+(2**8)* 70+  9, (2**17)*1+(2**8)* 88+ 77, 
(2**17)*0+(2**8)*  1+129, (2**17)*0+(2**8)* 20+ 76, (2**17)*0+(2**8)* 45+148, (2**17)*1+(2**8)* 85+ 58, 
(2**17)*0+(2**8)* 14+  5, (2**17)*0+(2**8)* 60+141, (2**17)*0+(2**8)* 74+  7, (2**17)*1+(2**8)* 82+ 62, 
(2**17)*0+(2**8)* 26+162, (2**17)*0+(2**8)* 95+123, (2**17)*0+(2**8)*100+138, (2**17)*1+(2**8)*115+134, 
(2**17)*0+(2**8)* 21+ 97, (2**17)*0+(2**8)* 56+  4, (2**17)*0+(2**8)* 75+ 23, (2**17)*1+(2**8)* 92+ 41, 
(2**17)*0+(2**8)*  7+119, (2**17)*0+(2**8)* 17+ 37, (2**17)*0+(2**8)* 35+ 83, (2**17)*1+(2**8)* 61+ 52, 
(2**17)*0+(2**8)* 17+147, (2**17)*0+(2**8)* 40+162, (2**17)*0+(2**8)* 86+101, (2**17)*1+(2**8)* 88+ 54, 
(2**17)*0+(2**8)*  4+121, (2**17)*0+(2**8)* 87+ 89, (2**17)*0+(2**8)*101+159, (2**17)*1+(2**8)*111+ 21, 
(2**17)*0+(2**8)* 15+ 84, (2**17)*0+(2**8)* 17+171, (2**17)*0+(2**8)* 93+162, (2**17)*1+(2**8)*119+166, 
(2**17)*0+(2**8)* 20+142, (2**17)*0+(2**8)* 44+ 60, (2**17)*0+(2**8)* 77+129, (2**17)*1+(2**8)* 86+174, 
(2**17)*0+(2**8)* 21+114, (2**17)*0+(2**8)* 85+ 99, (2**17)*0+(2**8)* 93+ 14, (2**17)*1+(2**8)*126+ 29, 
(2**17)*0+(2**8)*  7+  5, (2**17)*0+(2**8)* 22+154, (2**17)*0+(2**8)* 62+132, (2**17)*1+(2**8)* 73+ 61, 
(2**17)*0+(2**8)*  3+148, (2**17)*0+(2**8)* 22+121, (2**17)*0+(2**8)*106+147, (2**17)*1+(2**8)*136+109, 
(2**17)*0+(2**8)*  5+ 36, (2**17)*0+(2**8)*  9+ 81, (2**17)*0+(2**8)* 63+ 41, (2**17)*1+(2**8)* 73+ 93, 
(2**17)*0+(2**8)*  2+148, (2**17)*0+(2**8)*  7+ 25, (2**17)*0+(2**8)* 15+127, (2**17)*1+(2**8)*113+  1, 
(2**17)*0+(2**8)* 32+131, (2**17)*0+(2**8)* 72+ 23, (2**17)*0+(2**8)* 72+ 88, (2**17)*1+(2**8)*143+142, 
(2**17)*0+(2**8)* 17+121, (2**17)*0+(2**8)* 23+ 86, (2**17)*0+(2**8)* 91+ 64, (2**17)*1+(2**8)*117+ 33, 
(2**17)*0+(2**8)* 11+177, (2**17)*0+(2**8)* 40+ 68, (2**17)*0+(2**8)* 78+156, (2**17)*1+(2**8)*100+107, 
(2**17)*0+(2**8)*  1+ 63, (2**17)*0+(2**8)* 12+155, (2**17)*0+(2**8)* 23+106, (2**17)*1+(2**8)*121+149, 
(2**17)*0+(2**8)*  5+ 94, (2**17)*0+(2**8)* 16+131, (2**17)*0+(2**8)* 71+ 68, (2**17)*1+(2**8)* 85+166, 
(2**17)*0+(2**8)*  4+100, (2**17)*0+(2**8)*  5+ 51, (2**17)*0+(2**8)* 86+ 10, (2**17)*1+(2**8)*138+157, 
(2**17)*0+(2**8)* 10+114, (2**17)*0+(2**8)* 17+124, (2**17)*0+(2**8)* 89+ 27, (2**17)*1+(2**8)*116+ 75, 
(2**17)*0+(2**8)* 32+ 30, (2**17)*0+(2**8)* 61+158, (2**17)*0+(2**8)* 81+156, (2**17)*1+(2**8)* 96+ 80, 
(2**17)*0+(2**8)*  8+111, (2**17)*0+(2**8)* 12+ 67, (2**17)*0+(2**8)* 20+ 88, (2**17)*1+(2**8)*118+ 44, 
(2**17)*0+(2**8)*  2+ 48, (2**17)*0+(2**8)* 19+109, (2**17)*0+(2**8)* 82+  4, (2**17)*1+(2**8)*115+140, 
(2**17)*0+(2**8)* 67+ 49, (2**17)*0+(2**8)* 83+ 72, (2**17)*0+(2**8)* 90+113, (2**17)*1+(2**8)* 93+115, 
(2**17)*0+(2**8)* 84+ 31, (2**17)*0+(2**8)* 87+ 83, (2**17)*0+(2**8)* 89+ 54, (2**17)*1+(2**8)*114+ 80, 
(2**17)*0+(2**8)* 46+101, (2**17)*0+(2**8)* 72+ 67, (2**17)*0+(2**8)* 74+112, (2**17)*1+(2**8)* 93+ 19, 
(2**17)*0+(2**8)*  0+ 68, (2**17)*0+(2**8)*  8+154, (2**17)*0+(2**8)* 60+102, (2**17)*1+(2**8)* 79+164, 
(2**17)*0+(2**8)* 14+118, (2**17)*0+(2**8)* 26+144, (2**17)*0+(2**8)* 27+154, (2**17)*1+(2**8)* 47+108, 
(2**17)*0+(2**8)* 14+101, (2**17)*0+(2**8)* 94+132, (2**17)*0+(2**8)* 95+177, (2**17)*1+(2**8)*129+ 61, 
(2**17)*0+(2**8)* 15+122, (2**17)*0+(2**8)* 59+ 48, (2**17)*0+(2**8)* 89+119, (2**17)*1+(2**8)* 93+ 93, 
(2**17)*0+(2**8)*  4+ 59, (2**17)*0+(2**8)* 59+  5, (2**17)*0+(2**8)* 80+162, (2**17)*1+(2**8)* 95+114, 
(2**17)*0+(2**8)*  7+ 80, (2**17)*0+(2**8)* 81+103, (2**17)*0+(2**8)* 93+ 56, (2**17)*1+(2**8)*135+ 98, 
(2**17)*0+(2**8)*  6+167, (2**17)*0+(2**8)* 80+107, (2**17)*0+(2**8)* 83+163, (2**17)*1+(2**8)*140+ 61, 
(2**17)*0+(2**8)*  1+157, (2**17)*0+(2**8)* 13+138, (2**17)*0+(2**8)* 77+ 83, (2**17)*1+(2**8)*131+  7, 
(2**17)*0+(2**8)* 14+143, (2**17)*0+(2**8)* 22+  6, (2**17)*0+(2**8)* 48+ 86, (2**17)*1+(2**8)* 79+149, 
(2**17)*0+(2**8)*  2+ 53, (2**17)*0+(2**8)* 12+ 97, (2**17)*0+(2**8)* 88+ 26, (2**17)*1+(2**8)*128+ 35, 
(2**17)*0+(2**8)* 10+ 46, (2**17)*0+(2**8)* 72+  2, (2**17)*0+(2**8)* 81+127, (2**17)*1+(2**8)*137+ 92, 
(2**17)*0+(2**8)* 75+ 33, (2**17)*0+(2**8)* 76+ 37, (2**17)*0+(2**8)* 77+121, (2**17)*1+(2**8)*121+127, 
(2**17)*0+(2**8)* 88+ 79, (2**17)*0+(2**8)* 91+ 63, (2**17)*0+(2**8)* 96+ 88, (2**17)*1+(2**8)*128+ 49, 
(2**17)*0+(2**8)*  4+106, (2**17)*0+(2**8)*  8+ 70, (2**17)*0+(2**8)* 19+ 51, (2**17)*1+(2**8)* 53+132, 
(2**17)*0+(2**8)* 16+ 28, (2**17)*0+(2**8)* 22+142, (2**17)*0+(2**8)* 73+137, (2**17)*1+(2**8)*111+117, 
(2**17)*0+(2**8)*  6+166, (2**17)*0+(2**8)* 34+ 37, (2**17)*0+(2**8)* 50+139, (2**17)*1+(2**8)* 80+ 80, 
(2**17)*0+(2**8)*  1+ 76, (2**17)*0+(2**8)*  4+149, (2**17)*0+(2**8)* 64+164, (2**17)*1+(2**8)* 95+ 12, 
(2**17)*0+(2**8)*  6+ 85, (2**17)*0+(2**8)* 18+164, (2**17)*0+(2**8)* 51+129, (2**17)*1+(2**8)* 75+ 88, 
(2**17)*0+(2**8)*  6+ 71, (2**17)*0+(2**8)* 83+ 90, (2**17)*0+(2**8)* 99+177, (2**17)*1+(2**8)*125+ 91, 
(2**17)*0+(2**8)*  9+ 16, (2**17)*0+(2**8)* 15+ 31, (2**17)*0+(2**8)* 18+ 51, (2**17)*1+(2**8)*110+ 67, 
(2**17)*0+(2**8)*  9+126, (2**17)*0+(2**8)* 17+ 72, (2**17)*0+(2**8)* 31+104, (2**17)*1+(2**8)*141+144, 
(2**17)*0+(2**8)* 72+ 77, (2**17)*0+(2**8)* 82+ 96, (2**17)*0+(2**8)* 87+156, (2**17)*1+(2**8)*129+124, 
(2**17)*0+(2**8)* 21+113, (2**17)*0+(2**8)* 78+ 56, (2**17)*0+(2**8)* 85+ 50, (2**17)*1+(2**8)*139+131, 
(2**17)*0+(2**8)* 15+165, (2**17)*0+(2**8)* 17+ 43, (2**17)*0+(2**8)* 48+132, (2**17)*1+(2**8)* 81+ 14, 
(2**17)*0+(2**8)*  2+ 42, (2**17)*0+(2**8)* 33+135, (2**17)*0+(2**8)* 65+ 53, (2**17)*1+(2**8)* 83+ 63, 
(2**17)*0+(2**8)*  8+ 77, (2**17)*0+(2**8)* 62+ 61, (2**17)*0+(2**8)* 84+101, (2**17)*1+(2**8)* 85+172, 
(2**17)*0+(2**8)* 11+ 71, (2**17)*0+(2**8)* 13+ 86, (2**17)*0+(2**8)* 76+ 50, (2**17)*1+(2**8)*109+ 39, 
(2**17)*0+(2**8)* 16+ 69, (2**17)*0+(2**8)* 22+ 60, (2**17)*0+(2**8)* 50+146, (2**17)*1+(2**8)* 79+ 51, 
(2**17)*0+(2**8)* 19+ 90, (2**17)*0+(2**8)* 50+130, (2**17)*0+(2**8)* 76+155, (2**17)*1+(2**8)* 77+ 68, 
(2**17)*0+(2**8)* 18+ 52, (2**17)*0+(2**8)* 58+169, (2**17)*0+(2**8)* 72+ 87, (2**17)*1+(2**8)* 85+131, 
(2**17)*0+(2**8)* 18+127, (2**17)*0+(2**8)* 83+ 56, (2**17)*0+(2**8)* 97+147, (2**17)*1+(2**8)*140+101, 
(2**17)*0+(2**8)* 15+ 80, (2**17)*0+(2**8)* 79+139, (2**17)*0+(2**8)* 88+179, (2**17)*1+(2**8)*141+ 20, 
(2**17)*0+(2**8)* 11+ 15, (2**17)*0+(2**8)* 13+ 11, (2**17)*0+(2**8)* 74+115, (2**17)*1+(2**8)*109+120, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)* 32+  4, (2**17)*0+(2**8)* 58+ 73, (2**17)*1+(2**8)* 95+159, 
(2**17)*0+(2**8)*  6+ 32, (2**17)*0+(2**8)* 14+158, (2**17)*0+(2**8)* 68+ 97, (2**17)*1+(2**8)* 91+ 24, 
(2**17)*0+(2**8)*  0+133, (2**17)*0+(2**8)* 21+172, (2**17)*0+(2**8)* 74+143, (2**17)*1+(2**8)*113+ 36, 
(2**17)*0+(2**8)*  3+ 33, (2**17)*0+(2**8)* 11+159, (2**17)*0+(2**8)* 20+157, (2**17)*1+(2**8)* 37+ 61, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*0+(2**8)* 52+ 61, (2**17)*0+(2**8)* 73+ 62, (2**17)*1+(2**8)* 95+ 42, 
(2**17)*0+(2**8)*  3+100, (2**17)*0+(2**8)* 13+ 21, (2**17)*0+(2**8)* 34+ 93, (2**17)*1+(2**8)* 44+  9, 
(2**17)*0+(2**8)*  9+140, (2**17)*0+(2**8)* 84+172, (2**17)*0+(2**8)* 99+115, (2**17)*1+(2**8)*141+ 22, 
(2**17)*0+(2**8)* 18+ 32, (2**17)*0+(2**8)* 22+ 64, (2**17)*0+(2**8)* 62+163, (2**17)*1+(2**8)* 89+122, 
(2**17)*0+(2**8)* 78+  7, (2**17)*0+(2**8)* 81+ 21, (2**17)*0+(2**8)* 85+ 33, (2**17)*1+(2**8)*110+ 91, 
(2**17)*0+(2**8)* 80+104, (2**17)*0+(2**8)* 90+175, (2**17)*0+(2**8)* 91+ 84, (2**17)*1+(2**8)*129+ 48, 
(2**17)*0+(2**8)*  7+ 38, (2**17)*0+(2**8)* 80+ 24, (2**17)*0+(2**8)* 97+ 56, (2**17)*1+(2**8)*124+ 58, 
(2**17)*0+(2**8)* 12+109, (2**17)*0+(2**8)* 16+162, (2**17)*0+(2**8)* 64+ 80, (2**17)*1+(2**8)* 94+166, 
(2**17)*0+(2**8)*  2+106, (2**17)*0+(2**8)* 74+ 69, (2**17)*0+(2**8)* 82+145, (2**17)*1+(2**8)*119+156, 
(2**17)*0+(2**8)*  9+100, (2**17)*0+(2**8)* 12+ 34, (2**17)*0+(2**8)* 35+123, (2**17)*1+(2**8)*123+ 39, 
(2**17)*0+(2**8)* 11+ 17, (2**17)*0+(2**8)* 41+  5, (2**17)*0+(2**8)* 77+145, (2**17)*1+(2**8)*105+ 92, 
(2**17)*0+(2**8)* 14+142, (2**17)*0+(2**8)* 46+179, (2**17)*0+(2**8)* 83+ 70, (2**17)*1+(2**8)* 92+106, 
(2**17)*0+(2**8)*  6+ 18, (2**17)*0+(2**8)* 23+ 99, (2**17)*0+(2**8)* 76+ 49, (2**17)*1+(2**8)*112+118, 
(2**17)*0+(2**8)* 18+159, (2**17)*0+(2**8)* 22+176, (2**17)*0+(2**8)* 66+155, (2**17)*1+(2**8)* 91+ 55, 
(2**17)*0+(2**8)* 19+ 34, (2**17)*0+(2**8)* 45+ 90, (2**17)*0+(2**8)* 76+170, (2**17)*1+(2**8)* 77+ 46, 
(2**17)*0+(2**8)*  5+164, (2**17)*0+(2**8)* 16+166, (2**17)*0+(2**8)* 29+167, (2**17)*1+(2**8)* 51+ 70, 
(2**17)*0+(2**8)*  3+ 57, (2**17)*0+(2**8)* 12+ 61, (2**17)*0+(2**8)* 16+ 64, (2**17)*1+(2**8)*130+ 99, 
(2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 36+137, (2**17)*0+(2**8)* 73+ 92, (2**17)*1+(2**8)* 80+ 95, 
(2**17)*0+(2**8)* 16+168, (2**17)*0+(2**8)* 42+142, (2**17)*0+(2**8)* 76+ 72, (2**17)*1+(2**8)*105+ 16, 
(2**17)*0+(2**8)*  7+121, (2**17)*0+(2**8)* 19+ 50, (2**17)*0+(2**8)*107+168, (2**17)*1+(2**8)*121+105, 
(2**17)*0+(2**8)*  1+ 61, (2**17)*0+(2**8)* 19+164, (2**17)*0+(2**8)* 42+ 24, (2**17)*1+(2**8)* 80+  3, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)* 54+ 20, (2**17)*0+(2**8)* 83+109, (2**17)*1+(2**8)* 95+ 27, 
(2**17)*0+(2**8)*  2+ 82, (2**17)*0+(2**8)* 21+118, (2**17)*0+(2**8)* 90+ 82, (2**17)*1+(2**8)*127+ 55, 
(2**17)*0+(2**8)*  1+ 77, (2**17)*0+(2**8)*  8+ 24, (2**17)*0+(2**8)* 20+121, (2**17)*1+(2**8)*115+125, 
(2**17)*0+(2**8)* 31+ 67, (2**17)*0+(2**8)* 53+ 11, (2**17)*0+(2**8)* 84+119, (2**17)*1+(2**8)* 84+ 46, 
(2**17)*0+(2**8)* 18+ 36, (2**17)*0+(2**8)* 29+ 48, (2**17)*0+(2**8)* 48+ 83, (2**17)*1+(2**8)*102+ 33, 
(2**17)*0+(2**8)*  3+114, (2**17)*0+(2**8)* 87+126, (2**17)*0+(2**8)* 96+126, (2**17)*1+(2**8)*110+170, 
(2**17)*0+(2**8)* 21+ 66, (2**17)*0+(2**8)* 31+176, (2**17)*0+(2**8)* 70+ 25, (2**17)*1+(2**8)* 94+150, 
(2**17)*0+(2**8)* 10+ 31, (2**17)*0+(2**8)* 13+ 26, (2**17)*0+(2**8)* 86+ 77, (2**17)*1+(2**8)*142+ 22, 
(2**17)*0+(2**8)* 18+174, (2**17)*0+(2**8)* 75+ 83, (2**17)*0+(2**8)* 84+131, (2**17)*1+(2**8)*143+ 78, 
(2**17)*0+(2**8)*  2+ 51, (2**17)*0+(2**8)* 61+ 23, (2**17)*0+(2**8)* 79+ 13, (2**17)*1+(2**8)* 79+172, 
(2**17)*0+(2**8)* 22+ 39, (2**17)*0+(2**8)* 63+  6, (2**17)*0+(2**8)* 82+ 12, (2**17)*1+(2**8)* 91+143, 
(2**17)*0+(2**8)* 20+ 30, (2**17)*0+(2**8)* 20+108, (2**17)*0+(2**8)* 23+151, (2**17)*1+(2**8)* 39+ 33, 
(2**17)*0+(2**8)*  5+147, (2**17)*0+(2**8)* 10+117, (2**17)*0+(2**8)* 67+ 92, (2**17)*1+(2**8)* 72+  4, 
(2**17)*0+(2**8)* 20+172, (2**17)*0+(2**8)* 52+ 68, (2**17)*0+(2**8)* 73+ 28, (2**17)*1+(2**8)* 92+ 29, 
(2**17)*0+(2**8)* 10+126, (2**17)*0+(2**8)* 78+ 65, (2**17)*0+(2**8)* 90+100, (2**17)*1+(2**8)*137+153, 
(2**17)*0+(2**8)* 14+152, (2**17)*0+(2**8)* 15+ 75, (2**17)*0+(2**8)* 60+168, (2**17)*1+(2**8)* 82+ 32, 
(2**17)*0+(2**8)* 17+133, (2**17)*0+(2**8)* 28+175, (2**17)*0+(2**8)* 92+ 93, (2**17)*1+(2**8)*138+ 36, 
(2**17)*0+(2**8)*  9+ 25, (2**17)*0+(2**8)* 36+ 62, (2**17)*0+(2**8)* 76+ 91, (2**17)*1+(2**8)* 98+ 56, 
(2**17)*0+(2**8)*  6+ 58, (2**17)*0+(2**8)* 10+ 50, (2**17)*0+(2**8)* 55+ 38, (2**17)*1+(2**8)* 95+126, 
(2**17)*0+(2**8)* 15+106, (2**17)*0+(2**8)* 75+150, (2**17)*0+(2**8)* 78+169, (2**17)*1+(2**8)*127+131, 
(2**17)*0+(2**8)* 30+163, (2**17)*0+(2**8)* 36+ 34, (2**17)*0+(2**8)* 75+ 62, (2**17)*1+(2**8)* 86+ 98, 
(2**17)*0+(2**8)* 54+121, (2**17)*0+(2**8)* 77+154, (2**17)*0+(2**8)* 81+ 40, (2**17)*1+(2**8)* 97+119, 
(2**17)*0+(2**8)* 16+ 76, (2**17)*0+(2**8)* 72+145, (2**17)*0+(2**8)* 94+ 99, (2**17)*1+(2**8)*142+  9, 
(2**17)*0+(2**8)* 13+ 57, (2**17)*0+(2**8)* 73+129, (2**17)*0+(2**8)* 92+ 76, (2**17)*1+(2**8)*117+148, 
(2**17)*0+(2**8)*  2+  6, (2**17)*0+(2**8)* 10+ 61, (2**17)*0+(2**8)* 86+  5, (2**17)*1+(2**8)*132+141, 
(2**17)*0+(2**8)* 23+122, (2**17)*0+(2**8)* 28+137, (2**17)*0+(2**8)* 43+133, (2**17)*1+(2**8)* 98+162, 
(2**17)*0+(2**8)*  3+ 22, (2**17)*0+(2**8)* 20+ 40, (2**17)*0+(2**8)* 93+ 97, (2**17)*1+(2**8)*128+  4, 
(2**17)*0+(2**8)* 79+119, (2**17)*0+(2**8)* 89+ 37, (2**17)*0+(2**8)*107+ 83, (2**17)*1+(2**8)*133+ 52, 
(2**17)*0+(2**8)* 14+100, (2**17)*0+(2**8)* 16+ 53, (2**17)*0+(2**8)* 89+147, (2**17)*1+(2**8)*112+162, 
(2**17)*0+(2**8)* 15+ 88, (2**17)*0+(2**8)* 29+158, (2**17)*0+(2**8)* 39+ 20, (2**17)*1+(2**8)* 76+121, 
(2**17)*0+(2**8)* 21+161, (2**17)*0+(2**8)* 47+165, (2**17)*0+(2**8)* 87+ 84, (2**17)*1+(2**8)* 89+171, 
(2**17)*0+(2**8)*  5+128, (2**17)*0+(2**8)* 14+173, (2**17)*0+(2**8)* 92+142, (2**17)*1+(2**8)*116+ 60, 
(2**17)*0+(2**8)* 13+ 98, (2**17)*0+(2**8)* 21+ 13, (2**17)*0+(2**8)* 54+ 28, (2**17)*1+(2**8)* 93+114, 
(2**17)*0+(2**8)*  1+ 60, (2**17)*0+(2**8)* 79+  5, (2**17)*0+(2**8)* 94+154, (2**17)*1+(2**8)*134+132, 
(2**17)*0+(2**8)* 34+146, (2**17)*0+(2**8)* 64+108, (2**17)*0+(2**8)* 75+148, (2**17)*1+(2**8)* 94+121, 
(2**17)*0+(2**8)*  1+ 92, (2**17)*0+(2**8)* 77+ 36, (2**17)*0+(2**8)* 81+ 81, (2**17)*1+(2**8)*135+ 41, 
(2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 74+148, (2**17)*0+(2**8)* 79+ 25, (2**17)*1+(2**8)* 87+127, 


(2**17)*0+(2**8)* 26+150, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)*117+130, (2**17)*0+(2**8)*120+ 34, (2**17)*1+(2**8)*164+ 91, 
(2**17)*0+(2**8)* 10+ 25, (2**17)*0+(2**8)* 20+143, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 41+ 77, (2**17)*1+(2**8)*100+ 31, 
(2**17)*0+(2**8)* 16+  7, (2**17)*0+(2**8)* 27+159, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 51+ 69, (2**17)*1+(2**8)* 94+ 16, 
(2**17)*0+(2**8)*  2+131, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 68+176, (2**17)*0+(2**8)* 96+ 35, (2**17)*1+(2**8)*106+134, 
(2**17)*0+(2**8)* 33+ 18, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 82+139, (2**17)*0+(2**8)* 99+159, (2**17)*1+(2**8)*114+120, 
(2**17)*0+(2**8)*  3+ 76, (2**17)*0+(2**8)* 13+127, (2**17)*0+(2**8)* 24+ 68, (2**17)*0+(2**8)* 41+  0, (2**17)*1+(2**8)*120+105, 
(2**17)*0+(2**8)* 14+143, (2**17)*0+(2**8)* 32+118, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 76+169, (2**17)*1+(2**8)*111+ 52, 
(2**17)*0+(2**8)*  4+ 63, (2**17)*0+(2**8)* 28+ 22, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 89+107, (2**17)*1+(2**8)*124+133, 
(2**17)*0+(2**8)* 16+166, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)*108+  8, (2**17)*0+(2**8)*120+149, (2**17)*1+(2**8)*177+ 25, 
(2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 58+148, (2**17)*0+(2**8)*111+171, (2**17)*0+(2**8)*114+171, (2**17)*1+(2**8)*169+177, 
(2**17)*0+(2**8)*  1+ 14, (2**17)*0+(2**8)*  4+ 70, (2**17)*0+(2**8)*  5+ 88, (2**17)*0+(2**8)* 46+  0, (2**17)*1+(2**8)*127+  1, 
(2**17)*0+(2**8)* 19+100, (2**17)*0+(2**8)* 32+ 85, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 98+139, (2**17)*1+(2**8)*110+ 67, 
(2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)*105+167, (2**17)*0+(2**8)*116+ 40, (2**17)*0+(2**8)*123+ 91, (2**17)*1+(2**8)*168+ 99, 
(2**17)*0+(2**8)*  8+ 50, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)*106+ 73, (2**17)*0+(2**8)*136+158, (2**17)*1+(2**8)*156+116, 
(2**17)*0+(2**8)*  0+ 14, (2**17)*0+(2**8)* 18+113, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 63+ 50, (2**17)*1+(2**8)*157+ 66, 
(2**17)*0+(2**8)* 13+ 83, (2**17)*0+(2**8)* 30+ 92, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)*113+168, (2**17)*1+(2**8)*153+150, 
(2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 59+ 62, (2**17)*0+(2**8)* 96+ 68, (2**17)*0+(2**8)*101+120, (2**17)*1+(2**8)*163+ 43, 
(2**17)*0+(2**8)* 27+ 27, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 56+151, (2**17)*0+(2**8)* 98+ 87, (2**17)*1+(2**8)*139+ 61, 
(2**17)*0+(2**8)* 14+ 55, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)*113+ 26, (2**17)*0+(2**8)*115+137, (2**17)*1+(2**8)*171+ 81, 
(2**17)*0+(2**8)*  2+ 96, (2**17)*0+(2**8)* 28+ 80, (2**17)*0+(2**8)* 38+ 57, (2**17)*0+(2**8)* 55+  0, (2**17)*1+(2**8)*105+ 70, 
(2**17)*0+(2**8)* 11+ 25, (2**17)*0+(2**8)* 19+ 17, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 74+ 47, (2**17)*1+(2**8)*121+147, 
(2**17)*0+(2**8)*  0+153, (2**17)*0+(2**8)* 11+ 94, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 67+140, (2**17)*1+(2**8)* 98+ 12, 
(2**17)*0+(2**8)* 31+153, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 71+145, (2**17)*0+(2**8)*109+ 45, (2**17)*1+(2**8)*175+ 28, 
(2**17)*0+(2**8)*  9+ 22, (2**17)*0+(2**8)* 19+ 85, (2**17)*0+(2**8)* 45+ 92, (2**17)*0+(2**8)* 59+  0, (2**17)*1+(2**8)* 93+104, 
(2**17)*0+(2**8)* 35+102, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 94+ 18, (2**17)*0+(2**8)*107+ 37, (2**17)*1+(2**8)*142+ 49, 
(2**17)*0+(2**8)* 27+114, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 78+ 38, (2**17)*0+(2**8)*109+  2, (2**17)*1+(2**8)*114+145, 
(2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 92+145, (2**17)*0+(2**8)*119+ 59, (2**17)*0+(2**8)*142+ 43, (2**17)*1+(2**8)*173+122, 
(2**17)*0+(2**8)*  7+ 65, (2**17)*0+(2**8)* 13+ 84, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)*124+ 35, (2**17)*1+(2**8)*156+ 10, 
(2**17)*0+(2**8)* 25+166, (2**17)*0+(2**8)* 32+  5, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)*108+137, (2**17)*1+(2**8)*135+ 62, 
(2**17)*0+(2**8)*  5+119, (2**17)*0+(2**8)*  6+119, (2**17)*0+(2**8)* 14+ 37, (2**17)*0+(2**8)* 65+  0, (2**17)*1+(2**8)*125+ 71, 
(2**17)*0+(2**8)* 20+ 63, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 86+ 15, (2**17)*0+(2**8)*112+ 31, (2**17)*1+(2**8)*137+ 78, 
(2**17)*0+(2**8)*  3+ 64, (2**17)*0+(2**8)*  4+163, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)*136+ 93, (2**17)*1+(2**8)*170+117, 
(2**17)*0+(2**8)*  6+101, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)*107+165, (2**17)*0+(2**8)*115+ 95, (2**17)*1+(2**8)*154+107, 
(2**17)*0+(2**8)* 40+ 23, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)*105+ 56, (2**17)*0+(2**8)*106+ 44, (2**17)*1+(2**8)*125+147, 
(2**17)*0+(2**8)* 12+144, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 88+162, (2**17)*0+(2**8)*101+ 24, (2**17)*1+(2**8)*167+ 86, 
(2**17)*0+(2**8)* 22+ 76, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)*104+115, (2**17)*0+(2**8)*118+ 87, (2**17)*1+(2**8)*126+139, 
(2**17)*0+(2**8)* 51+148, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 95+ 18, (2**17)*0+(2**8)*111+115, (2**17)*1+(2**8)*115+139, 
(2**17)*0+(2**8)*  4+ 72, (2**17)*0+(2**8)* 61+ 98, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)*100+143, (2**17)*1+(2**8)*121+ 35, 
(2**17)*0+(2**8)* 10+ 82, (2**17)*0+(2**8)* 50+ 21, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 97+ 52, (2**17)*1+(2**8)*127+ 22, 
(2**17)*0+(2**8)* 26+166, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)*110+ 51, (2**17)*0+(2**8)*138+179, (2**17)*1+(2**8)*145+ 48, 
(2**17)*0+(2**8)* 20+ 44, (2**17)*0+(2**8)* 70+ 68, (2**17)*0+(2**8)* 75+ 56, (2**17)*0+(2**8)* 76+  0, (2**17)*1+(2**8)*105+169, 
(2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)*107+175, (2**17)*0+(2**8)*121+138, (2**17)*0+(2**8)*147+ 84, (2**17)*1+(2**8)*148+ 34, 
(2**17)*0+(2**8)* 20+119, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)*106+156, (2**17)*0+(2**8)*117+123, (2**17)*1+(2**8)*176+ 37, 
(2**17)*0+(2**8)* 14+ 30, (2**17)*0+(2**8)* 21+ 25, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)*149+ 58, (2**17)*1+(2**8)*179+112, 
(2**17)*0+(2**8)*  8+ 30, (2**17)*0+(2**8)* 19+ 74, (2**17)*0+(2**8)* 39+  4, (2**17)*0+(2**8)* 80+  0, (2**17)*1+(2**8)*115+ 54, 
(2**17)*0+(2**8)*  5+ 34, (2**17)*0+(2**8)* 18+ 29, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)* 91+ 26, (2**17)*1+(2**8)*112+ 89, 
(2**17)*0+(2**8)* 71+ 36, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)* 97+ 33, (2**17)*0+(2**8)*111+165, (2**17)*1+(2**8)*123+ 13, 
(2**17)*0+(2**8)* 65+170, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 90+ 48, (2**17)*0+(2**8)*116+ 83, (2**17)*1+(2**8)*140+120, 
(2**17)*0+(2**8)* 14+102, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)* 90+ 52, (2**17)*0+(2**8)*100+ 90, (2**17)*1+(2**8)*125+106, 
(2**17)*0+(2**8)*  5+ 93, (2**17)*0+(2**8)* 33+148, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)* 90+ 57, (2**17)*1+(2**8)*119+ 10, 
(2**17)*0+(2**8)*  1+156, (2**17)*0+(2**8)* 11+124, (2**17)*0+(2**8)* 12+ 58, (2**17)*0+(2**8)* 60+ 74, (2**17)*1+(2**8)* 86+  0, 
(2**17)*0+(2**8)*  1+ 20, (2**17)*0+(2**8)*  3+ 32, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*111+122, (2**17)*1+(2**8)*175+115, 
(2**17)*0+(2**8)* 17+175, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)* 95+118, (2**17)*0+(2**8)*163+150, (2**17)*1+(2**8)*177+ 71, 
(2**17)*0+(2**8)* 10+123, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)*113+ 73, (2**17)*0+(2**8)*130+ 69, (2**17)*1+(2**8)*158+ 99, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  3+145, (2**17)*0+(2**8)*  6+ 46, (2**17)*0+(2**8)*  8+131, (2**17)*1+(2**8)* 83+ 25, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 88+  3, (2**17)*0+(2**8)*115+174, (2**17)*0+(2**8)*120+  3, (2**17)*1+(2**8)*143+ 83, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  6+172, (2**17)*0+(2**8)* 28+ 88, (2**17)*0+(2**8)* 30+ 16, (2**17)*1+(2**8)*132+  6, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)* 12+ 53, (2**17)*0+(2**8)* 26+154, (2**17)*0+(2**8)* 60+ 53, (2**17)*1+(2**8)* 93+ 86, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 29+ 28, (2**17)*0+(2**8)* 94+160, (2**17)*0+(2**8)*113+104, (2**17)*1+(2**8)*125+140, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 29+ 56, (2**17)*0+(2**8)* 54+ 87, (2**17)*0+(2**8)*107+ 53, (2**17)*1+(2**8)*134+ 45, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 38+  1, (2**17)*0+(2**8)* 57+150, (2**17)*0+(2**8)*102+180, (2**17)*1+(2**8)*111+156, 
(2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)* 12+171, (2**17)*0+(2**8)* 61+ 39, (2**17)*0+(2**8)*121+112, (2**17)*1+(2**8)*160+148, 
(2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 12+ 34, (2**17)*0+(2**8)* 12+ 15, (2**17)*0+(2**8)* 35+ 49, (2**17)*1+(2**8)*155+101, 
(2**17)*0+(2**8)*  1+ 40, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 29+162, (2**17)*0+(2**8)* 34+ 66, (2**17)*1+(2**8)* 91+ 17, 
(2**17)*0+(2**8)*  3+ 90, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 23+162, (2**17)*0+(2**8)*108+ 36, (2**17)*1+(2**8)*123+113, 
(2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 47+137, (2**17)*0+(2**8)* 72+145, (2**17)*0+(2**8)*103+107, (2**17)*1+(2**8)*107+ 52, 
(2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 15+ 26, (2**17)*0+(2**8)* 97+127, (2**17)*0+(2**8)*114+176, (2**17)*1+(2**8)*171+ 39, 
(2**17)*0+(2**8)*  9+123, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 34+116, (2**17)*0+(2**8)* 49+ 15, (2**17)*1+(2**8)*120+136, 
(2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 32+103, (2**17)*0+(2**8)* 43+ 29, (2**17)*0+(2**8)* 96+ 98, (2**17)*1+(2**8)*121+124, 
(2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 26+ 63, (2**17)*0+(2**8)* 79+ 69, (2**17)*0+(2**8)* 84+ 44, (2**17)*1+(2**8)*112+173, 
(2**17)*0+(2**8)*  1+132, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 20+  8, (2**17)*0+(2**8)*103+123, (2**17)*1+(2**8)*122+ 69, 
(2**17)*0+(2**8)*  2+137, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 17+ 82, (2**17)*0+(2**8)* 24+142, (2**17)*1+(2**8)* 28+ 31, 
(2**17)*0+(2**8)*  2+  4, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 53+112, (2**17)*0+(2**8)*124+ 87, (2**17)*1+(2**8)*129+134, 
(2**17)*0+(2**8)* 18+ 92, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 27+165, (2**17)*0+(2**8)* 35+ 39, (2**17)*1+(2**8)* 62+108, 
(2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 22+142, (2**17)*0+(2**8)* 75+ 65, (2**17)*0+(2**8)* 99+ 94, (2**17)*1+(2**8)* 99+153, 
(2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 23+176, (2**17)*0+(2**8)* 77+  7, (2**17)*0+(2**8)*112+109, (2**17)*1+(2**8)*159+ 52, 
(2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 26+121, (2**17)*0+(2**8)*104+102, (2**17)*0+(2**8)*119+145, (2**17)*1+(2**8)*144+137, 
(2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 24+128, (2**17)*0+(2**8)* 28+126, (2**17)*0+(2**8)* 97+ 63, (2**17)*1+(2**8)*126+ 81, 
(2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 41+ 88, (2**17)*0+(2**8)* 44+156, (2**17)*0+(2**8)*103+ 76, (2**17)*1+(2**8)*105+138, 
(2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 82+  5, (2**17)*0+(2**8)* 92+ 51, (2**17)*0+(2**8)*112+122, (2**17)*1+(2**8)*138+100, 
(2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 64+ 49, (2**17)*0+(2**8)* 80+178, (2**17)*0+(2**8)* 92+ 32, (2**17)*1+(2**8)*103+166, 
(2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 72+ 62, (2**17)*0+(2**8)*106+122, (2**17)*0+(2**8)*124+127, (2**17)*1+(2**8)*166+167, 
(2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 55+177, (2**17)*0+(2**8)* 90+ 80, (2**17)*0+(2**8)* 99+144, (2**17)*1+(2**8)*124+ 84, 
(2**17)*0+(2**8)* 27+  1, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 97+ 79, (2**17)*0+(2**8)*123+109, (2**17)*1+(2**8)*152+  8, 
(2**17)*0+(2**8)* 18+  3, (2**17)*0+(2**8)* 28+121, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)*101+ 95, (2**17)*1+(2**8)*159+165, 
(2**17)*0+(2**8)* 10+ 81, (2**17)*0+(2**8)* 29+167, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 33+ 33, (2**17)*1+(2**8)* 99+119, 
(2**17)*0+(2**8)*  8+166, (2**17)*0+(2**8)* 23+ 59, (2**17)*0+(2**8)* 31+168, (2**17)*0+(2**8)* 32+  0, (2**17)*1+(2**8)* 32+162, 
(2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 42+118, (2**17)*0+(2**8)*101+130, (2**17)*0+(2**8)*115+177, (2**17)*1+(2**8)*174+121, 
(2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 95+ 89, (2**17)*0+(2**8)* 97+  4, (2**17)*0+(2**8)*105+ 77, (2**17)*1+(2**8)*146+111, 
(2**17)*0+(2**8)*  0+149, (2**17)*0+(2**8)* 19+108, (2**17)*0+(2**8)* 32+179, (2**17)*0+(2**8)* 35+  0, (2**17)*1+(2**8)*133+ 81, 
(2**17)*0+(2**8)* 27+129, (2**17)*0+(2**8)* 30+ 33, (2**17)*0+(2**8)* 74+ 90, (2**17)*0+(2**8)*116+150, (2**17)*1+(2**8)*126+  0, 
(2**17)*0+(2**8)* 10+ 30, (2**17)*0+(2**8)*100+ 25, (2**17)*0+(2**8)*110+143, (2**17)*0+(2**8)*127+  0, (2**17)*1+(2**8)*131+ 77, 
(2**17)*0+(2**8)*  4+ 15, (2**17)*0+(2**8)*106+  7, (2**17)*0+(2**8)*117+159, (2**17)*0+(2**8)*128+  0, (2**17)*1+(2**8)*141+ 69, 
(2**17)*0+(2**8)*  6+ 34, (2**17)*0+(2**8)* 16+133, (2**17)*0+(2**8)* 92+131, (2**17)*0+(2**8)*129+  0, (2**17)*1+(2**8)*158+176, 
(2**17)*0+(2**8)*  9+158, (2**17)*0+(2**8)* 24+119, (2**17)*0+(2**8)*123+ 18, (2**17)*0+(2**8)*130+  0, (2**17)*1+(2**8)*172+139, 
(2**17)*0+(2**8)* 30+104, (2**17)*0+(2**8)* 93+ 76, (2**17)*0+(2**8)*103+127, (2**17)*0+(2**8)*114+ 68, (2**17)*1+(2**8)*131+  0, 
(2**17)*0+(2**8)* 21+ 51, (2**17)*0+(2**8)*104+143, (2**17)*0+(2**8)*122+118, (2**17)*0+(2**8)*132+  0, (2**17)*1+(2**8)*166+169, 
(2**17)*0+(2**8)* 34+132, (2**17)*0+(2**8)* 94+ 63, (2**17)*0+(2**8)*118+ 22, (2**17)*0+(2**8)*133+  0, (2**17)*1+(2**8)*179+107, 
(2**17)*0+(2**8)* 18+  7, (2**17)*0+(2**8)* 30+148, (2**17)*0+(2**8)* 87+ 24, (2**17)*0+(2**8)*106+166, (2**17)*1+(2**8)*134+  0, 
(2**17)*0+(2**8)* 21+170, (2**17)*0+(2**8)* 24+170, (2**17)*0+(2**8)* 79+176, (2**17)*0+(2**8)*135+  0, (2**17)*1+(2**8)*148+148, 
(2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 91+ 14, (2**17)*0+(2**8)* 94+ 70, (2**17)*0+(2**8)* 95+ 88, (2**17)*1+(2**8)*136+  0, 
(2**17)*0+(2**8)*  8+138, (2**17)*0+(2**8)* 20+ 66, (2**17)*0+(2**8)*109+100, (2**17)*0+(2**8)*122+ 85, (2**17)*1+(2**8)*137+  0, 
(2**17)*0+(2**8)* 15+166, (2**17)*0+(2**8)* 26+ 39, (2**17)*0+(2**8)* 33+ 90, (2**17)*0+(2**8)* 78+ 98, (2**17)*1+(2**8)*138+  0, 
(2**17)*0+(2**8)* 16+ 72, (2**17)*0+(2**8)* 46+157, (2**17)*0+(2**8)* 66+115, (2**17)*0+(2**8)* 98+ 50, (2**17)*1+(2**8)*139+  0, 
(2**17)*0+(2**8)* 67+ 65, (2**17)*0+(2**8)* 90+ 14, (2**17)*0+(2**8)*108+113, (2**17)*0+(2**8)*140+  0, (2**17)*1+(2**8)*153+ 50, 
(2**17)*0+(2**8)* 23+167, (2**17)*0+(2**8)* 63+149, (2**17)*0+(2**8)*103+ 83, (2**17)*0+(2**8)*120+ 92, (2**17)*1+(2**8)*141+  0, 
(2**17)*0+(2**8)*  6+ 67, (2**17)*0+(2**8)* 11+119, (2**17)*0+(2**8)* 73+ 42, (2**17)*0+(2**8)*142+  0, (2**17)*1+(2**8)*149+ 62, 
(2**17)*0+(2**8)*  8+ 86, (2**17)*0+(2**8)* 49+ 60, (2**17)*0+(2**8)*117+ 27, (2**17)*0+(2**8)*143+  0, (2**17)*1+(2**8)*146+151, 
(2**17)*0+(2**8)* 23+ 25, (2**17)*0+(2**8)* 25+136, (2**17)*0+(2**8)* 81+ 80, (2**17)*0+(2**8)*104+ 55, (2**17)*1+(2**8)*144+  0, 
(2**17)*0+(2**8)* 15+ 69, (2**17)*0+(2**8)* 92+ 96, (2**17)*0+(2**8)*118+ 80, (2**17)*0+(2**8)*128+ 57, (2**17)*1+(2**8)*145+  0, 
(2**17)*0+(2**8)* 31+146, (2**17)*0+(2**8)*101+ 25, (2**17)*0+(2**8)*109+ 17, (2**17)*0+(2**8)*146+  0, (2**17)*1+(2**8)*164+ 47, 
(2**17)*0+(2**8)*  8+ 11, (2**17)*0+(2**8)* 90+153, (2**17)*0+(2**8)*101+ 94, (2**17)*0+(2**8)*147+  0, (2**17)*1+(2**8)*157+140, 
(2**17)*0+(2**8)* 19+ 44, (2**17)*0+(2**8)* 85+ 27, (2**17)*0+(2**8)*121+153, (2**17)*0+(2**8)*148+  0, (2**17)*1+(2**8)*161+145, 
(2**17)*0+(2**8)*  3+103, (2**17)*0+(2**8)* 99+ 22, (2**17)*0+(2**8)*109+ 85, (2**17)*0+(2**8)*135+ 92, (2**17)*1+(2**8)*149+  0, 
(2**17)*0+(2**8)*  4+ 17, (2**17)*0+(2**8)* 17+ 36, (2**17)*0+(2**8)* 52+ 48, (2**17)*0+(2**8)*125+102, (2**17)*1+(2**8)*150+  0, 
(2**17)*0+(2**8)* 19+  1, (2**17)*0+(2**8)* 24+144, (2**17)*0+(2**8)*117+114, (2**17)*0+(2**8)*151+  0, (2**17)*1+(2**8)*168+ 38, 
(2**17)*0+(2**8)*  2+144, (2**17)*0+(2**8)* 29+ 58, (2**17)*0+(2**8)* 52+ 42, (2**17)*0+(2**8)* 83+121, (2**17)*1+(2**8)*152+  0, 
(2**17)*0+(2**8)* 34+ 34, (2**17)*0+(2**8)* 66+  9, (2**17)*0+(2**8)* 97+ 65, (2**17)*0+(2**8)*103+ 84, (2**17)*1+(2**8)*153+  0, 
(2**17)*0+(2**8)* 18+136, (2**17)*0+(2**8)* 45+ 61, (2**17)*0+(2**8)*115+166, (2**17)*0+(2**8)*122+  5, (2**17)*1+(2**8)*154+  0, 
(2**17)*0+(2**8)* 35+ 70, (2**17)*0+(2**8)* 95+119, (2**17)*0+(2**8)* 96+119, (2**17)*0+(2**8)*104+ 37, (2**17)*1+(2**8)*155+  0, 
(2**17)*0+(2**8)* 22+ 30, (2**17)*0+(2**8)* 47+ 77, (2**17)*0+(2**8)*110+ 63, (2**17)*0+(2**8)*156+  0, (2**17)*1+(2**8)*176+ 15, 
(2**17)*0+(2**8)* 46+ 92, (2**17)*0+(2**8)* 80+116, (2**17)*0+(2**8)* 93+ 64, (2**17)*0+(2**8)* 94+163, (2**17)*1+(2**8)*157+  0, 
(2**17)*0+(2**8)* 17+164, (2**17)*0+(2**8)* 25+ 94, (2**17)*0+(2**8)* 64+106, (2**17)*0+(2**8)* 96+101, (2**17)*1+(2**8)*158+  0, 
(2**17)*0+(2**8)* 15+ 55, (2**17)*0+(2**8)* 16+ 43, (2**17)*0+(2**8)* 35+146, (2**17)*0+(2**8)*130+ 23, (2**17)*1+(2**8)*159+  0, 
(2**17)*0+(2**8)* 11+ 23, (2**17)*0+(2**8)* 77+ 85, (2**17)*0+(2**8)*102+144, (2**17)*0+(2**8)*160+  0, (2**17)*1+(2**8)*178+162, 
(2**17)*0+(2**8)* 14+114, (2**17)*0+(2**8)* 28+ 86, (2**17)*0+(2**8)* 36+138, (2**17)*0+(2**8)*112+ 76, (2**17)*1+(2**8)*161+  0, 
(2**17)*0+(2**8)*  5+ 17, (2**17)*0+(2**8)* 21+114, (2**17)*0+(2**8)* 25+138, (2**17)*0+(2**8)*141+148, (2**17)*1+(2**8)*162+  0, 
(2**17)*0+(2**8)* 10+142, (2**17)*0+(2**8)* 31+ 34, (2**17)*0+(2**8)* 94+ 72, (2**17)*0+(2**8)*151+ 98, (2**17)*1+(2**8)*163+  0, 
(2**17)*0+(2**8)*  7+ 51, (2**17)*0+(2**8)* 37+ 21, (2**17)*0+(2**8)*100+ 82, (2**17)*0+(2**8)*140+ 21, (2**17)*1+(2**8)*164+  0, 
(2**17)*0+(2**8)* 20+ 50, (2**17)*0+(2**8)* 48+178, (2**17)*0+(2**8)* 55+ 47, (2**17)*0+(2**8)*116+166, (2**17)*1+(2**8)*165+  0, 
(2**17)*0+(2**8)* 15+168, (2**17)*0+(2**8)*110+ 44, (2**17)*0+(2**8)*160+ 68, (2**17)*0+(2**8)*165+ 56, (2**17)*1+(2**8)*166+  0, 
(2**17)*0+(2**8)* 17+174, (2**17)*0+(2**8)* 31+137, (2**17)*0+(2**8)* 57+ 83, (2**17)*0+(2**8)* 58+ 33, (2**17)*1+(2**8)*167+  0, 
(2**17)*0+(2**8)* 16+155, (2**17)*0+(2**8)* 27+122, (2**17)*0+(2**8)* 86+ 36, (2**17)*0+(2**8)*110+119, (2**17)*1+(2**8)*168+  0, 
(2**17)*0+(2**8)* 59+ 57, (2**17)*0+(2**8)* 89+111, (2**17)*0+(2**8)*104+ 30, (2**17)*0+(2**8)*111+ 25, (2**17)*1+(2**8)*169+  0, 
(2**17)*0+(2**8)* 25+ 53, (2**17)*0+(2**8)* 98+ 30, (2**17)*0+(2**8)*109+ 74, (2**17)*0+(2**8)*129+  4, (2**17)*1+(2**8)*170+  0, 
(2**17)*0+(2**8)*  1+ 25, (2**17)*0+(2**8)* 22+ 88, (2**17)*0+(2**8)* 95+ 34, (2**17)*0+(2**8)*108+ 29, (2**17)*1+(2**8)*171+  0, 
(2**17)*0+(2**8)*  7+ 32, (2**17)*0+(2**8)* 21+164, (2**17)*0+(2**8)* 33+ 12, (2**17)*0+(2**8)*161+ 36, (2**17)*1+(2**8)*172+  0, 
(2**17)*0+(2**8)*  0+ 47, (2**17)*0+(2**8)* 26+ 82, (2**17)*0+(2**8)* 50+119, (2**17)*0+(2**8)*155+170, (2**17)*1+(2**8)*173+  0, 
(2**17)*0+(2**8)*  0+ 51, (2**17)*0+(2**8)* 10+ 89, (2**17)*0+(2**8)* 35+105, (2**17)*0+(2**8)*104+102, (2**17)*1+(2**8)*174+  0, 
(2**17)*0+(2**8)*  0+ 56, (2**17)*0+(2**8)* 29+  9, (2**17)*0+(2**8)* 95+ 93, (2**17)*0+(2**8)*123+148, (2**17)*1+(2**8)*175+  0, 
(2**17)*0+(2**8)* 91+156, (2**17)*0+(2**8)*101+124, (2**17)*0+(2**8)*102+ 58, (2**17)*0+(2**8)*150+ 74, (2**17)*1+(2**8)*176+  0, 
(2**17)*0+(2**8)* 21+121, (2**17)*0+(2**8)* 85+114, (2**17)*0+(2**8)* 91+ 20, (2**17)*0+(2**8)* 93+ 32, (2**17)*1+(2**8)*177+  0, 
(2**17)*0+(2**8)*  5+117, (2**17)*0+(2**8)* 73+149, (2**17)*0+(2**8)* 87+ 70, (2**17)*0+(2**8)*107+175, (2**17)*1+(2**8)*178+  0, 
(2**17)*0+(2**8)* 23+ 72, (2**17)*0+(2**8)* 40+ 68, (2**17)*0+(2**8)* 68+ 98, (2**17)*0+(2**8)*100+123, (2**17)*1+(2**8)*179+  0, 
(2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)* 93+145, (2**17)*0+(2**8)* 96+ 46, (2**17)*0+(2**8)* 98+131, (2**17)*1+(2**8)*173+ 25, 
(2**17)*0+(2**8)* 25+173, (2**17)*0+(2**8)* 30+  2, (2**17)*0+(2**8)* 53+ 82, (2**17)*0+(2**8)* 91+  0, (2**17)*1+(2**8)*178+  3, 
(2**17)*0+(2**8)* 42+  5, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)* 96+172, (2**17)*0+(2**8)*118+ 88, (2**17)*1+(2**8)*120+ 16, 
(2**17)*0+(2**8)*  3+ 85, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*102+ 53, (2**17)*0+(2**8)*116+154, (2**17)*1+(2**8)*150+ 53, 
(2**17)*0+(2**8)*  4+159, (2**17)*0+(2**8)* 23+103, (2**17)*0+(2**8)* 35+139, (2**17)*0+(2**8)* 94+  0, (2**17)*1+(2**8)*119+ 28, 
(2**17)*0+(2**8)* 17+ 52, (2**17)*0+(2**8)* 44+ 44, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*119+ 56, (2**17)*1+(2**8)*144+ 87, 
(2**17)*0+(2**8)* 12+179, (2**17)*0+(2**8)* 21+155, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*128+  1, (2**17)*1+(2**8)*147+150, 
(2**17)*0+(2**8)* 31+111, (2**17)*0+(2**8)* 70+147, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*102+171, (2**17)*1+(2**8)*151+ 39, 
(2**17)*0+(2**8)* 65+100, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*102+ 34, (2**17)*0+(2**8)*102+ 15, (2**17)*1+(2**8)*125+ 49, 
(2**17)*0+(2**8)*  1+ 16, (2**17)*0+(2**8)* 91+ 40, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*119+162, (2**17)*1+(2**8)*124+ 66, 
(2**17)*0+(2**8)* 18+ 35, (2**17)*0+(2**8)* 33+112, (2**17)*0+(2**8)* 93+ 90, (2**17)*0+(2**8)*100+  0, (2**17)*1+(2**8)*113+162, 
(2**17)*0+(2**8)* 13+106, (2**17)*0+(2**8)* 17+ 51, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*137+137, (2**17)*1+(2**8)*162+145, 
(2**17)*0+(2**8)*  7+126, (2**17)*0+(2**8)* 24+175, (2**17)*0+(2**8)* 81+ 38, (2**17)*0+(2**8)*102+  0, (2**17)*1+(2**8)*105+ 26, 
(2**17)*0+(2**8)* 30+135, (2**17)*0+(2**8)* 99+123, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*124+116, (2**17)*1+(2**8)*139+ 15, 
(2**17)*0+(2**8)*  6+ 97, (2**17)*0+(2**8)* 31+123, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*122+103, (2**17)*1+(2**8)*133+ 29, 
(2**17)*0+(2**8)* 22+172, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*116+ 63, (2**17)*0+(2**8)*169+ 69, (2**17)*1+(2**8)*174+ 44, 
(2**17)*0+(2**8)* 13+122, (2**17)*0+(2**8)* 32+ 68, (2**17)*0+(2**8)* 91+132, (2**17)*0+(2**8)*106+  0, (2**17)*1+(2**8)*110+  8, 
(2**17)*0+(2**8)* 92+137, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*107+ 82, (2**17)*0+(2**8)*114+142, (2**17)*1+(2**8)*118+ 31, 
(2**17)*0+(2**8)* 34+ 86, (2**17)*0+(2**8)* 39+133, (2**17)*0+(2**8)* 92+  4, (2**17)*0+(2**8)*108+  0, (2**17)*1+(2**8)*143+112, 
(2**17)*0+(2**8)*108+ 92, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*117+165, (2**17)*0+(2**8)*125+ 39, (2**17)*1+(2**8)*152+108, 
(2**17)*0+(2**8)*  9+ 93, (2**17)*0+(2**8)*  9+152, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*112+142, (2**17)*1+(2**8)*165+ 65, 
(2**17)*0+(2**8)* 22+108, (2**17)*0+(2**8)* 69+ 51, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*113+176, (2**17)*1+(2**8)*167+  7, 
(2**17)*0+(2**8)* 14+101, (2**17)*0+(2**8)* 29+144, (2**17)*0+(2**8)* 54+136, (2**17)*0+(2**8)*112+  0, (2**17)*1+(2**8)*116+121, 
(2**17)*0+(2**8)*  7+ 62, (2**17)*0+(2**8)* 36+ 80, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*114+128, (2**17)*1+(2**8)*118+126, 
(2**17)*0+(2**8)* 13+ 75, (2**17)*0+(2**8)* 15+137, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*131+ 88, (2**17)*1+(2**8)*134+156, 
(2**17)*0+(2**8)*  2+ 50, (2**17)*0+(2**8)* 22+121, (2**17)*0+(2**8)* 48+ 99, (2**17)*0+(2**8)*115+  0, (2**17)*1+(2**8)*172+  5, 
(2**17)*0+(2**8)*  2+ 31, (2**17)*0+(2**8)* 13+165, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*154+ 49, (2**17)*1+(2**8)*170+178, 
(2**17)*0+(2**8)* 16+121, (2**17)*0+(2**8)* 34+126, (2**17)*0+(2**8)* 76+166, (2**17)*0+(2**8)*117+  0, (2**17)*1+(2**8)*162+ 62, 
(2**17)*0+(2**8)*  0+ 79, (2**17)*0+(2**8)*  9+143, (2**17)*0+(2**8)* 34+ 83, (2**17)*0+(2**8)*118+  0, (2**17)*1+(2**8)*145+177, 
(2**17)*0+(2**8)*  7+ 78, (2**17)*0+(2**8)* 33+108, (2**17)*0+(2**8)* 62+  7, (2**17)*0+(2**8)*117+  1, (2**17)*1+(2**8)*119+  0, 
(2**17)*0+(2**8)* 11+ 94, (2**17)*0+(2**8)* 69+164, (2**17)*0+(2**8)*108+  3, (2**17)*0+(2**8)*118+121, (2**17)*1+(2**8)*120+  0, 
(2**17)*0+(2**8)*  9+118, (2**17)*0+(2**8)*100+ 81, (2**17)*0+(2**8)*119+167, (2**17)*0+(2**8)*121+  0, (2**17)*1+(2**8)*123+ 33, 
(2**17)*0+(2**8)* 98+166, (2**17)*0+(2**8)*113+ 59, (2**17)*0+(2**8)*121+168, (2**17)*0+(2**8)*122+  0, (2**17)*1+(2**8)*122+162, 
(2**17)*0+(2**8)* 11+129, (2**17)*0+(2**8)* 25+176, (2**17)*0+(2**8)* 84+120, (2**17)*0+(2**8)*123+  0, (2**17)*1+(2**8)*132+118, 
(2**17)*0+(2**8)*  5+ 88, (2**17)*0+(2**8)*  7+  3, (2**17)*0+(2**8)* 15+ 76, (2**17)*0+(2**8)* 56+110, (2**17)*1+(2**8)*124+  0, 
(2**17)*0+(2**8)* 43+ 80, (2**17)*0+(2**8)* 90+149, (2**17)*0+(2**8)*109+108, (2**17)*0+(2**8)*122+179, (2**17)*1+(2**8)*125+  0, 


(2**17)*0+(2**8)* 15+100, (2**17)*0+(2**8)* 24+ 67, (2**17)*0+(2**8)* 33+ 57, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)*108+119, (2**17)*0+(2**8)*130+157, (2**17)*0+(2**8)*140+173, (2**17)*0+(2**8)*148+105, (2**17)*1+(2**8)*209+102, 
(2**17)*0+(2**8)*  7+ 69, (2**17)*0+(2**8)*  9+ 13, (2**17)*0+(2**8)* 11+131, (2**17)*0+(2**8)* 33+ 67, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 44+ 37, (2**17)*0+(2**8)* 97+173, (2**17)*0+(2**8)*108+ 78, (2**17)*1+(2**8)*132+ 34, 
(2**17)*0+(2**8)*  8+ 89, (2**17)*0+(2**8)* 14+ 26, (2**17)*0+(2**8)* 33+ 78, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 64+ 47, (2**17)*0+(2**8)*110+179, (2**17)*0+(2**8)*114+129, (2**17)*0+(2**8)*142+ 18, (2**17)*1+(2**8)*200+170, 
(2**17)*0+(2**8)* 17+ 93, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)*120+164, (2**17)*0+(2**8)*125+109, (2**17)*0+(2**8)*130+ 73, (2**17)*0+(2**8)*134+130, (2**17)*0+(2**8)*135+122, (2**17)*0+(2**8)*165+180, (2**17)*1+(2**8)*212+106, 
(2**17)*0+(2**8)* 18+ 25, (2**17)*0+(2**8)* 25+ 17, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 96+179, (2**17)*0+(2**8)*115+177, (2**17)*0+(2**8)*119+ 63, (2**17)*0+(2**8)*122+ 70, (2**17)*0+(2**8)*126+ 61, (2**17)*1+(2**8)*163+ 12, 
(2**17)*0+(2**8)* 24+105, (2**17)*0+(2**8)* 25+ 80, (2**17)*0+(2**8)* 31+ 60, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)*130+105, (2**17)*0+(2**8)*136+  6, (2**17)*0+(2**8)*137+ 27, (2**17)*0+(2**8)*156+101, (2**17)*1+(2**8)*202+ 69, 
(2**17)*0+(2**8)* 10+ 90, (2**17)*0+(2**8)* 12+ 50, (2**17)*0+(2**8)* 17+176, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 50+ 92, (2**17)*0+(2**8)*114+ 43, (2**17)*0+(2**8)*128+123, (2**17)*0+(2**8)*133+143, (2**17)*1+(2**8)*206+171, 
(2**17)*0+(2**8)* 10+ 31, (2**17)*0+(2**8)* 18+114, (2**17)*0+(2**8)* 25+ 92, (2**17)*0+(2**8)* 27+149, (2**17)*0+(2**8)* 30+ 43, (2**17)*0+(2**8)* 31+ 22, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)*153+130, (2**17)*1+(2**8)*205+144, 
(2**17)*0+(2**8)*  3+177, (2**17)*0+(2**8)*  8+ 44, (2**17)*0+(2**8)*  8+ 49, (2**17)*0+(2**8)* 22+ 28, (2**17)*0+(2**8)* 35+123, (2**17)*0+(2**8)* 38+ 65, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)*116+ 61, (2**17)*1+(2**8)*187+179, 
(2**17)*0+(2**8)*  0+ 39, (2**17)*0+(2**8)* 22+ 33, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 67+ 32, (2**17)*0+(2**8)* 77+171, (2**17)*0+(2**8)*115+ 59, (2**17)*0+(2**8)*119+ 79, (2**17)*0+(2**8)*138+165, (2**17)*1+(2**8)*139+ 85, 
(2**17)*0+(2**8)*  1+ 29, (2**17)*0+(2**8)* 24+117, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)*121+ 31, (2**17)*0+(2**8)*125+ 41, (2**17)*0+(2**8)*131+ 94, (2**17)*0+(2**8)*138+ 66, (2**17)*0+(2**8)*159+134, (2**17)*1+(2**8)*211+  7, 
(2**17)*0+(2**8)*  4+ 53, (2**17)*0+(2**8)*  9+150, (2**17)*0+(2**8)* 11+ 46, (2**17)*0+(2**8)* 11+ 68, (2**17)*0+(2**8)* 15+168, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 82+144, (2**17)*0+(2**8)*124+122, (2**17)*1+(2**8)*164+ 31, 
(2**17)*0+(2**8)*  5+ 37, (2**17)*0+(2**8)* 11+101, (2**17)*0+(2**8)* 13+ 81, (2**17)*0+(2**8)* 25+140, (2**17)*0+(2**8)* 33+173, (2**17)*0+(2**8)* 41+128, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 94+ 57, (2**17)*1+(2**8)*143+ 52, 
(2**17)*0+(2**8)* 31+ 20, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 81+  7, (2**17)*0+(2**8)*111+ 48, (2**17)*0+(2**8)*111+111, (2**17)*0+(2**8)*115+ 26, (2**17)*0+(2**8)*123+160, (2**17)*0+(2**8)*142+ 82, (2**17)*1+(2**8)*144+130, 
(2**17)*0+(2**8)* 17+166, (2**17)*0+(2**8)* 28+159, (2**17)*0+(2**8)* 29+176, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 69+ 14, (2**17)*0+(2**8)* 89+ 48, (2**17)*0+(2**8)*115+ 33, (2**17)*0+(2**8)*121+143, (2**17)*1+(2**8)*123+ 56, 
(2**17)*0+(2**8)* 23+153, (2**17)*0+(2**8)* 27+113, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)*112+101, (2**17)*0+(2**8)*123+ 53, (2**17)*0+(2**8)*139+ 72, (2**17)*0+(2**8)*140+ 59, (2**17)*0+(2**8)*168+112, (2**17)*1+(2**8)*188+ 84, 
(2**17)*0+(2**8)* 13+123, (2**17)*0+(2**8)* 19+128, (2**17)*0+(2**8)* 27+131, (2**17)*0+(2**8)* 29+ 35, (2**17)*0+(2**8)* 41+171, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)*117+161, (2**17)*0+(2**8)*123+ 36, (2**17)*1+(2**8)*210+ 26, 
(2**17)*0+(2**8)*  2+ 15, (2**17)*0+(2**8)*  5+176, (2**17)*0+(2**8)* 26+102, (2**17)*0+(2**8)* 35+ 44, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 60+150, (2**17)*0+(2**8)* 90+ 43, (2**17)*0+(2**8)*131+  3, (2**17)*1+(2**8)*137+160, 
(2**17)*0+(2**8)*  4+121, (2**17)*0+(2**8)* 14+ 20, (2**17)*0+(2**8)* 20+ 42, (2**17)*0+(2**8)* 23+168, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 58+158, (2**17)*0+(2**8)* 99+ 86, (2**17)*0+(2**8)*109+113, (2**17)*1+(2**8)*122+ 65, 
(2**17)*0+(2**8)*  2+ 94, (2**17)*0+(2**8)*  5+ 39, (2**17)*0+(2**8)*  7+178, (2**17)*0+(2**8)*  9+ 52, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 59+ 98, (2**17)*0+(2**8)*135+ 21, (2**17)*0+(2**8)*139+ 26, (2**17)*1+(2**8)*199+ 97, 
(2**17)*0+(2**8)* 10+145, (2**17)*0+(2**8)* 19+ 61, (2**17)*0+(2**8)* 23+ 83, (2**17)*0+(2**8)* 32+152, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 63+ 56, (2**17)*0+(2**8)*110+ 61, (2**17)*0+(2**8)*119+154, (2**17)*1+(2**8)*200+ 92, 
(2**17)*0+(2**8)*  3+115, (2**17)*0+(2**8)*  4+168, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 62+  4, (2**17)*0+(2**8)*110+134, (2**17)*0+(2**8)*114+ 38, (2**17)*0+(2**8)*123+ 91, (2**17)*0+(2**8)*126+114, (2**17)*1+(2**8)*183+ 36, 
(2**17)*0+(2**8)*  3+151, (2**17)*0+(2**8)* 17+ 29, (2**17)*0+(2**8)* 21+115, (2**17)*0+(2**8)* 29+132, (2**17)*0+(2**8)* 49+  5, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)*102+118, (2**17)*0+(2**8)*134+106, (2**17)*1+(2**8)*134+ 71, 
(2**17)*0+(2**8)*  1+118, (2**17)*0+(2**8)* 27+ 55, (2**17)*0+(2**8)* 42+133, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 79+152, (2**17)*0+(2**8)*117+143, (2**17)*0+(2**8)*127+145, (2**17)*0+(2**8)*135+ 29, (2**17)*1+(2**8)*135+ 39, 
(2**17)*0+(2**8)*  1+178, (2**17)*0+(2**8)*  6+ 62, (2**17)*0+(2**8)* 20+ 31, (2**17)*0+(2**8)* 21+169, (2**17)*0+(2**8)* 30+153, (2**17)*0+(2**8)* 35+ 17, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 86+ 45, (2**17)*1+(2**8)*170+139, 
(2**17)*0+(2**8)*  1+139, (2**17)*0+(2**8)*  1+120, (2**17)*0+(2**8)* 11+ 88, (2**17)*0+(2**8)* 32+142, (2**17)*0+(2**8)* 51+ 92, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)*125+104, (2**17)*0+(2**8)*133+ 25, (2**17)*1+(2**8)*184+158, 
(2**17)*0+(2**8)* 16+ 24, (2**17)*0+(2**8)* 17+106, (2**17)*0+(2**8)* 28+142, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 76+ 48, (2**17)*0+(2**8)*108+ 22, (2**17)*0+(2**8)*122+138, (2**17)*0+(2**8)*143+ 11, (2**17)*1+(2**8)*160+147, 
(2**17)*0+(2**8)* 35+ 25, (2**17)*0+(2**8)* 43+ 76, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)*108+  1, (2**17)*0+(2**8)*114+ 91, (2**17)*0+(2**8)*118+104, (2**17)*0+(2**8)*124+ 91, (2**17)*0+(2**8)*140+ 26, (2**17)*1+(2**8)*191+106, 
(2**17)*0+(2**8)*  2+ 38, (2**17)*0+(2**8)* 10+ 32, (2**17)*0+(2**8)* 30+157, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)*118+ 86, (2**17)*0+(2**8)*126+ 67, (2**17)*0+(2**8)*140+127, (2**17)*0+(2**8)*155+ 51, (2**17)*1+(2**8)*180+174, 
(2**17)*0+(2**8)*  5+140, (2**17)*0+(2**8)* 10+114, (2**17)*0+(2**8)* 27+ 47, (2**17)*0+(2**8)* 30+114, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 75+147, (2**17)*0+(2**8)*110+159, (2**17)*0+(2**8)*119+156, (2**17)*1+(2**8)*167+ 75, 
(2**17)*0+(2**8)* 53+158, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)*108+156, (2**17)*0+(2**8)*116+121, (2**17)*0+(2**8)*116+ 37, (2**17)*0+(2**8)*121+102, (2**17)*0+(2**8)*130+177, (2**17)*0+(2**8)*137+165, (2**17)*1+(2**8)*207+ 26, 
(2**17)*0+(2**8)*  1+174, (2**17)*0+(2**8)*  4+ 77, (2**17)*0+(2**8)* 10+ 64, (2**17)*0+(2**8)* 33+ 75, (2**17)*0+(2**8)* 52+ 42, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)*134+140, (2**17)*0+(2**8)*140+ 38, (2**17)*1+(2**8)*193+100, 
(2**17)*0+(2**8)*  6+145, (2**17)*0+(2**8)* 23+ 71, (2**17)*0+(2**8)* 66+ 94, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 88+ 61, (2**17)*0+(2**8)*115+ 99, (2**17)*0+(2**8)*129+ 10, (2**17)*0+(2**8)*130+ 68, (2**17)*1+(2**8)*140+112, 
(2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 83+ 78, (2**17)*0+(2**8)*110+ 77, (2**17)*0+(2**8)*111+164, (2**17)*0+(2**8)*116+ 97, (2**17)*0+(2**8)*122+167, (2**17)*0+(2**8)*124+171, (2**17)*0+(2**8)*138+168, (2**17)*1+(2**8)*146+ 75, 
(2**17)*0+(2**8)*  3+ 36, (2**17)*0+(2**8)*  6+ 47, (2**17)*0+(2**8)* 19+ 92, (2**17)*0+(2**8)* 23+119, (2**17)*0+(2**8)* 23+ 41, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)*108+ 81, (2**17)*0+(2**8)*151+132, (2**17)*1+(2**8)*208+ 58, 
(2**17)*0+(2**8)*  0+  1, (2**17)*0+(2**8)*  3+ 87, (2**17)*0+(2**8)*  3+ 80, (2**17)*0+(2**8)* 13+ 82, (2**17)*0+(2**8)* 27+162, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)*132+166, (2**17)*0+(2**8)*144+129, (2**17)*1+(2**8)*204+121, 
(2**17)*0+(2**8)*  5+ 45, (2**17)*0+(2**8)* 13+  5, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)*109+  6, (2**17)*0+(2**8)*112+  8, (2**17)*0+(2**8)*132+ 21, (2**17)*0+(2**8)*134+147, (2**17)*0+(2**8)*155+154, (2**17)*1+(2**8)*214+ 25, 
(2**17)*0+(2**8)*  5+104, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)*109+ 81, (2**17)*0+(2**8)*124+ 52, (2**17)*0+(2**8)*125+168, (2**17)*0+(2**8)*127+120, (2**17)*0+(2**8)*132+ 51, (2**17)*0+(2**8)*173+ 30, (2**17)*1+(2**8)*211+138, 
(2**17)*0+(2**8)* 25+162, (2**17)*0+(2**8)* 34+133, (2**17)*0+(2**8)* 35+ 96, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 74+ 34, (2**17)*0+(2**8)*117+160, (2**17)*0+(2**8)*119+127, (2**17)*0+(2**8)*120+139, (2**17)*1+(2**8)*152+139, 
(2**17)*0+(2**8)* 20+114, (2**17)*0+(2**8)* 42+144, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)*123+ 52, (2**17)*0+(2**8)*128+152, (2**17)*0+(2**8)*130+ 60, (2**17)*0+(2**8)*137+ 62, (2**17)*0+(2**8)*138+ 28, (2**17)*1+(2**8)*194+ 17, 
(2**17)*0+(2**8)* 20+177, (2**17)*0+(2**8)* 26+ 49, (2**17)*0+(2**8)* 58+151, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)*104+ 84, (2**17)*0+(2**8)*119+ 54, (2**17)*0+(2**8)*123+  8, (2**17)*0+(2**8)*128+107, (2**17)*1+(2**8)*133+ 11, 
(2**17)*0+(2**8)*  9+ 20, (2**17)*0+(2**8)* 30+ 36, (2**17)*0+(2**8)* 34+173, (2**17)*0+(2**8)* 49+ 77, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)*112+115, (2**17)*0+(2**8)*133+134, (2**17)*0+(2**8)*133+171, (2**17)*1+(2**8)*201+ 94, 
(2**17)*0+(2**8)*  0+ 20, (2**17)*0+(2**8)* 10+ 12, (2**17)*0+(2**8)* 29+ 69, (2**17)*0+(2**8)* 31+144, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)*110+ 79, (2**17)*0+(2**8)*130+164, (2**17)*0+(2**8)*148+ 93, (2**17)*1+(2**8)*189+169, 
(2**17)*0+(2**8)*  4+ 98, (2**17)*0+(2**8)* 12+  8, (2**17)*0+(2**8)* 18+ 56, (2**17)*0+(2**8)* 34+ 78, (2**17)*0+(2**8)* 34+ 16, (2**17)*0+(2**8)* 69+136, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)* 88+100, (2**17)*1+(2**8)*132+ 91, 
(2**17)*0+(2**8)*  8+149, (2**17)*0+(2**8)* 15+175, (2**17)*0+(2**8)* 64+ 66, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)* 82+ 97, (2**17)*0+(2**8)*116+ 28, (2**17)*0+(2**8)*120+ 87, (2**17)*0+(2**8)*128+100, (2**17)*1+(2**8)*134+137, 
(2**17)*0+(2**8)*  2+ 21, (2**17)*0+(2**8)*  9+ 39, (2**17)*0+(2**8)* 33+ 59, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)*106+ 20, (2**17)*0+(2**8)*126+172, (2**17)*0+(2**8)*138+ 54, (2**17)*0+(2**8)*138+156, (2**17)*1+(2**8)*163+135, 
(2**17)*0+(2**8)*  8+172, (2**17)*0+(2**8)*  8+ 15, (2**17)*0+(2**8)* 24+ 91, (2**17)*0+(2**8)* 24+166, (2**17)*0+(2**8)* 77+ 52, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)*141+ 45, (2**17)*0+(2**8)*142+ 50, (2**17)*1+(2**8)*173+122, 
(2**17)*0+(2**8)* 13+ 25, (2**17)*0+(2**8)* 21+162, (2**17)*0+(2**8)* 26+ 39, (2**17)*0+(2**8)* 54+137, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 91+ 28, (2**17)*0+(2**8)*115+ 63, (2**17)*0+(2**8)*134+131, (2**17)*1+(2**8)*143+ 20, 
(2**17)*0+(2**8)* 12+131, (2**17)*0+(2**8)* 13+159, (2**17)*0+(2**8)* 21+177, (2**17)*0+(2**8)* 27+155, (2**17)*0+(2**8)* 71+120, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)*112+146, (2**17)*0+(2**8)*129+ 90, (2**17)*1+(2**8)*180+ 97, 
(2**17)*0+(2**8)*  3+154, (2**17)*0+(2**8)*  9+137, (2**17)*0+(2**8)* 20+ 12, (2**17)*0+(2**8)* 28+ 28, (2**17)*0+(2**8)* 56+ 25, (2**17)*0+(2**8)* 73+156, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*121+ 90, (2**17)*1+(2**8)*131+124, 
(2**17)*0+(2**8)* 20+126, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)*113+ 66, (2**17)*0+(2**8)*115+117, (2**17)*0+(2**8)*122+  6, (2**17)*0+(2**8)*137+164, (2**17)*0+(2**8)*140+ 69, (2**17)*0+(2**8)*145+ 21, (2**17)*1+(2**8)*215+ 24, 
(2**17)*0+(2**8)*  1+156, (2**17)*0+(2**8)* 12+139, (2**17)*0+(2**8)* 33+132, (2**17)*0+(2**8)* 34+172, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*122+ 35, (2**17)*0+(2**8)*131+ 38, (2**17)*0+(2**8)*165+ 93, (2**17)*1+(2**8)*192+108, 
(2**17)*0+(2**8)*  7+ 38, (2**17)*0+(2**8)* 14+ 61, (2**17)*0+(2**8)* 21+ 28, (2**17)*0+(2**8)* 39+ 54, (2**17)*0+(2**8)* 87+173, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)*129+ 59, (2**17)*0+(2**8)*131+112, (2**17)*1+(2**8)*141+ 73, 
(2**17)*0+(2**8)*  7+165, (2**17)*0+(2**8)*  9+156, (2**17)*0+(2**8)* 13+ 57, (2**17)*0+(2**8)* 28+ 34, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)*108+139, (2**17)*0+(2**8)*117+ 17, (2**17)*0+(2**8)*169+ 26, (2**17)*1+(2**8)*186+ 89, 
(2**17)*0+(2**8)* 16+ 64, (2**17)*0+(2**8)* 68+161, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)*124+115, (2**17)*0+(2**8)*124+102, (2**17)*0+(2**8)*125+ 26, (2**17)*0+(2**8)*127+176, (2**17)*0+(2**8)*140+ 18, (2**17)*1+(2**8)*213+ 54, 
(2**17)*0+(2**8)* 18+115, (2**17)*0+(2**8)* 31+ 82, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)*101+139, (2**17)*0+(2**8)*109+ 45, (2**17)*0+(2**8)*120+146, (2**17)*0+(2**8)*135+ 56, (2**17)*0+(2**8)*137+ 92, (2**17)*1+(2**8)*171+ 40, 
(2**17)*0+(2**8)* 16+ 25, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*105+158, (2**17)*0+(2**8)*123+ 33, (2**17)*0+(2**8)*126+173, (2**17)*0+(2**8)*126+180, (2**17)*0+(2**8)*130+  1, (2**17)*0+(2**8)*130+ 13, (2**17)*1+(2**8)*176+ 81, 
(2**17)*0+(2**8)*  9+132, (2**17)*0+(2**8)* 34+ 50, (2**17)*0+(2**8)* 61+ 44, (2**17)*0+(2**8)* 85+ 65, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*110+120, (2**17)*0+(2**8)*120+ 43, (2**17)*0+(2**8)*124+110, (2**17)*1+(2**8)*127+ 26, 
(2**17)*0+(2**8)*  0+ 71, (2**17)*0+(2**8)*  5+  7, (2**17)*0+(2**8)* 25+122, (2**17)*0+(2**8)* 28+ 50, (2**17)*0+(2**8)* 31+ 55, (2**17)*0+(2**8)* 34+ 20, (2**17)*0+(2**8)* 67+ 12, (2**17)*0+(2**8)* 94+  0, (2**17)*1+(2**8)*203+ 11, 
(2**17)*0+(2**8)*  3+176, (2**17)*0+(2**8)*  4+ 74, (2**17)*0+(2**8)* 12+166, (2**17)*0+(2**8)* 19+ 35, (2**17)*0+(2**8)* 39+ 85, (2**17)*0+(2**8)* 74+ 87, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*113+ 99, (2**17)*1+(2**8)*124+165, 
(2**17)*0+(2**8)*  6+154, (2**17)*0+(2**8)* 25+125, (2**17)*0+(2**8)* 33+ 79, (2**17)*0+(2**8)* 35+104, (2**17)*0+(2**8)* 71+ 95, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*110+100, (2**17)*0+(2**8)*136+ 49, (2**17)*1+(2**8)*188+  8, 
(2**17)*0+(2**8)* 18+141, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*100+  9, (2**17)*0+(2**8)*111+137, (2**17)*0+(2**8)*113+116, (2**17)*0+(2**8)*122+169, (2**17)*0+(2**8)*128+ 87, (2**17)*0+(2**8)*129+155, (2**17)*1+(2**8)*158+ 96, 
(2**17)*0+(2**8)*  0+ 57, (2**17)*0+(2**8)* 12+ 30, (2**17)*0+(2**8)* 29+148, (2**17)*0+(2**8)* 30+ 92, (2**17)*0+(2**8)* 32+ 78, (2**17)*0+(2**8)* 84+ 32, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*141+114, (2**17)*1+(2**8)*145+ 73, 
(2**17)*0+(2**8)*  4+ 39, (2**17)*0+(2**8)* 22+174, (2**17)*0+(2**8)* 32+158, (2**17)*0+(2**8)* 73+ 46, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*109+157, (2**17)*0+(2**8)*136+170, (2**17)*0+(2**8)*139+179, (2**17)*1+(2**8)*174+157, 
(2**17)*0+(2**8)* 10+ 76, (2**17)*0+(2**8)* 45+ 78, (2**17)*0+(2**8)* 78+169, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*114+ 48, (2**17)*0+(2**8)*116+115, (2**17)*0+(2**8)*131+147, (2**17)*0+(2**8)*142+113, (2**17)*1+(2**8)*143+161, 
(2**17)*0+(2**8)* 26+ 97, (2**17)*0+(2**8)* 31+118, (2**17)*0+(2**8)* 35+ 41, (2**17)*0+(2**8)* 70+ 94, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*115+137, (2**17)*0+(2**8)*122+ 77, (2**17)*0+(2**8)*125+118, (2**17)*1+(2**8)*215+ 54, 
(2**17)*0+(2**8)* 20+121, (2**17)*0+(2**8)* 21+ 44, (2**17)*0+(2**8)* 24+170, (2**17)*0+(2**8)* 29+ 98, (2**17)*0+(2**8)* 70+ 93, (2**17)*0+(2**8)* 87+171, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*113+ 10, (2**17)*1+(2**8)*127+171, 
(2**17)*0+(2**8)* 46+143, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*114+109, (2**17)*0+(2**8)*114+150, (2**17)*0+(2**8)*118+ 19, (2**17)*0+(2**8)*136+ 74, (2**17)*0+(2**8)*141+ 40, (2**17)*0+(2**8)*142+ 88, (2**17)*1+(2**8)*197+  9, 
(2**17)*0+(2**8)*  4+108, (2**17)*0+(2**8)*  6+  3, (2**17)*0+(2**8)* 53+ 40, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*113+ 60, (2**17)*0+(2**8)*122+ 56, (2**17)*0+(2**8)*125+158, (2**17)*0+(2**8)*134+ 87, (2**17)*1+(2**8)*203+ 42, 
(2**17)*0+(2**8)* 12+172, (2**17)*0+(2**8)* 18+ 93, (2**17)*0+(2**8)* 19+142, (2**17)*0+(2**8)* 28+ 99, (2**17)*0+(2**8)* 93+ 42, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*119+177, (2**17)*0+(2**8)*143+  4, (2**17)*1+(2**8)*156+153, 
(2**17)*0+(2**8)* 13+ 77, (2**17)*0+(2**8)* 19+ 68, (2**17)*0+(2**8)* 24+137, (2**17)*0+(2**8)* 28+  7, (2**17)*0+(2**8)* 46+104, (2**17)*0+(2**8)* 90+144, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*124+156, (2**17)*1+(2**8)*136+ 30, 
(2**17)*0+(2**8)* 10+  5, (2**17)*0+(2**8)* 15+ 38, (2**17)*0+(2**8)* 19+ 98, (2**17)*0+(2**8)* 21+ 56, (2**17)*0+(2**8)* 54+ 29, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*129+145, (2**17)*0+(2**8)*139+171, (2**17)*1+(2**8)*206+143, 
(2**17)*0+(2**8)*  0+118, (2**17)*0+(2**8)* 22+156, (2**17)*0+(2**8)* 32+172, (2**17)*0+(2**8)* 40+104, (2**17)*0+(2**8)*101+101, (2**17)*0+(2**8)*123+100, (2**17)*0+(2**8)*132+ 67, (2**17)*0+(2**8)*141+ 57, (2**17)*1+(2**8)*144+  0, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*0+(2**8)* 24+ 33, (2**17)*0+(2**8)*115+ 69, (2**17)*0+(2**8)*117+ 13, (2**17)*0+(2**8)*119+131, (2**17)*0+(2**8)*141+ 67, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*152+ 37, (2**17)*1+(2**8)*205+173, 
(2**17)*0+(2**8)*  2+178, (2**17)*0+(2**8)*  6+128, (2**17)*0+(2**8)* 34+ 17, (2**17)*0+(2**8)* 92+169, (2**17)*0+(2**8)*116+ 89, (2**17)*0+(2**8)*122+ 26, (2**17)*0+(2**8)*141+ 78, (2**17)*0+(2**8)*146+  0, (2**17)*1+(2**8)*172+ 47, 
(2**17)*0+(2**8)* 12+163, (2**17)*0+(2**8)* 17+108, (2**17)*0+(2**8)* 22+ 72, (2**17)*0+(2**8)* 26+129, (2**17)*0+(2**8)* 27+121, (2**17)*0+(2**8)* 57+179, (2**17)*0+(2**8)*104+105, (2**17)*0+(2**8)*125+ 93, (2**17)*1+(2**8)*147+  0, 
(2**17)*0+(2**8)*  7+176, (2**17)*0+(2**8)* 11+ 62, (2**17)*0+(2**8)* 14+ 69, (2**17)*0+(2**8)* 18+ 60, (2**17)*0+(2**8)* 55+ 11, (2**17)*0+(2**8)*126+ 25, (2**17)*0+(2**8)*133+ 17, (2**17)*0+(2**8)*148+  0, (2**17)*1+(2**8)*204+179, 
(2**17)*0+(2**8)* 22+104, (2**17)*0+(2**8)* 28+  5, (2**17)*0+(2**8)* 29+ 26, (2**17)*0+(2**8)* 48+100, (2**17)*0+(2**8)* 94+ 68, (2**17)*0+(2**8)*132+105, (2**17)*0+(2**8)*133+ 80, (2**17)*0+(2**8)*139+ 60, (2**17)*1+(2**8)*149+  0, 
(2**17)*0+(2**8)*  6+ 42, (2**17)*0+(2**8)* 20+122, (2**17)*0+(2**8)* 25+142, (2**17)*0+(2**8)* 98+170, (2**17)*0+(2**8)*118+ 90, (2**17)*0+(2**8)*120+ 50, (2**17)*0+(2**8)*125+176, (2**17)*0+(2**8)*150+  0, (2**17)*1+(2**8)*158+ 92, 
(2**17)*0+(2**8)* 45+129, (2**17)*0+(2**8)* 97+143, (2**17)*0+(2**8)*118+ 31, (2**17)*0+(2**8)*126+114, (2**17)*0+(2**8)*133+ 92, (2**17)*0+(2**8)*135+149, (2**17)*0+(2**8)*138+ 43, (2**17)*0+(2**8)*139+ 22, (2**17)*1+(2**8)*151+  0, 
(2**17)*0+(2**8)*  8+ 60, (2**17)*0+(2**8)* 79+178, (2**17)*0+(2**8)*111+177, (2**17)*0+(2**8)*116+ 44, (2**17)*0+(2**8)*116+ 49, (2**17)*0+(2**8)*130+ 28, (2**17)*0+(2**8)*143+123, (2**17)*0+(2**8)*146+ 65, (2**17)*1+(2**8)*152+  0, 
(2**17)*0+(2**8)*  7+ 58, (2**17)*0+(2**8)* 11+ 78, (2**17)*0+(2**8)* 30+164, (2**17)*0+(2**8)* 31+ 84, (2**17)*0+(2**8)*108+ 39, (2**17)*0+(2**8)*130+ 33, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*175+ 32, (2**17)*1+(2**8)*185+171, 
(2**17)*0+(2**8)* 13+ 30, (2**17)*0+(2**8)* 17+ 40, (2**17)*0+(2**8)* 23+ 93, (2**17)*0+(2**8)* 30+ 65, (2**17)*0+(2**8)* 51+133, (2**17)*0+(2**8)*103+  6, (2**17)*0+(2**8)*109+ 29, (2**17)*0+(2**8)*132+117, (2**17)*1+(2**8)*154+  0, 
(2**17)*0+(2**8)* 16+121, (2**17)*0+(2**8)* 56+ 30, (2**17)*0+(2**8)*112+ 53, (2**17)*0+(2**8)*117+150, (2**17)*0+(2**8)*119+ 46, (2**17)*0+(2**8)*119+ 68, (2**17)*0+(2**8)*123+168, (2**17)*0+(2**8)*155+  0, (2**17)*1+(2**8)*190+144, 
(2**17)*0+(2**8)* 35+ 51, (2**17)*0+(2**8)*113+ 37, (2**17)*0+(2**8)*119+101, (2**17)*0+(2**8)*121+ 81, (2**17)*0+(2**8)*133+140, (2**17)*0+(2**8)*141+173, (2**17)*0+(2**8)*149+128, (2**17)*0+(2**8)*156+  0, (2**17)*1+(2**8)*202+ 57, 
(2**17)*0+(2**8)*  3+ 47, (2**17)*0+(2**8)*  3+110, (2**17)*0+(2**8)*  7+ 25, (2**17)*0+(2**8)* 15+159, (2**17)*0+(2**8)* 34+ 81, (2**17)*0+(2**8)* 36+129, (2**17)*0+(2**8)*139+ 20, (2**17)*0+(2**8)*157+  0, (2**17)*1+(2**8)*189+  7, 
(2**17)*0+(2**8)*  7+ 32, (2**17)*0+(2**8)* 13+142, (2**17)*0+(2**8)* 15+ 55, (2**17)*0+(2**8)*125+166, (2**17)*0+(2**8)*136+159, (2**17)*0+(2**8)*137+176, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*177+ 14, (2**17)*1+(2**8)*197+ 48, 
(2**17)*0+(2**8)*  4+100, (2**17)*0+(2**8)* 15+ 52, (2**17)*0+(2**8)* 31+ 71, (2**17)*0+(2**8)* 32+ 58, (2**17)*0+(2**8)* 60+111, (2**17)*0+(2**8)* 80+ 83, (2**17)*0+(2**8)*131+153, (2**17)*0+(2**8)*135+113, (2**17)*1+(2**8)*159+  0, 
(2**17)*0+(2**8)*  9+160, (2**17)*0+(2**8)* 15+ 35, (2**17)*0+(2**8)*102+ 25, (2**17)*0+(2**8)*121+123, (2**17)*0+(2**8)*127+128, (2**17)*0+(2**8)*135+131, (2**17)*0+(2**8)*137+ 35, (2**17)*0+(2**8)*149+171, (2**17)*1+(2**8)*160+  0, 
(2**17)*0+(2**8)* 23+  2, (2**17)*0+(2**8)* 29+159, (2**17)*0+(2**8)*110+ 15, (2**17)*0+(2**8)*113+176, (2**17)*0+(2**8)*134+102, (2**17)*0+(2**8)*143+ 44, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*168+150, (2**17)*1+(2**8)*198+ 43, 
(2**17)*0+(2**8)*  1+112, (2**17)*0+(2**8)* 14+ 64, (2**17)*0+(2**8)*112+121, (2**17)*0+(2**8)*122+ 20, (2**17)*0+(2**8)*128+ 42, (2**17)*0+(2**8)*131+168, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*166+158, (2**17)*1+(2**8)*207+ 86, 
(2**17)*0+(2**8)* 27+ 20, (2**17)*0+(2**8)* 31+ 25, (2**17)*0+(2**8)* 91+ 96, (2**17)*0+(2**8)*110+ 94, (2**17)*0+(2**8)*113+ 39, (2**17)*0+(2**8)*115+178, (2**17)*0+(2**8)*117+ 52, (2**17)*0+(2**8)*163+  0, (2**17)*1+(2**8)*167+ 98, 
(2**17)*0+(2**8)*  2+ 60, (2**17)*0+(2**8)* 11+153, (2**17)*0+(2**8)* 92+ 91, (2**17)*0+(2**8)*118+145, (2**17)*0+(2**8)*127+ 61, (2**17)*0+(2**8)*131+ 83, (2**17)*0+(2**8)*140+152, (2**17)*0+(2**8)*164+  0, (2**17)*1+(2**8)*171+ 56, 
(2**17)*0+(2**8)*  2+133, (2**17)*0+(2**8)*  6+ 37, (2**17)*0+(2**8)* 15+ 90, (2**17)*0+(2**8)* 18+113, (2**17)*0+(2**8)* 75+ 35, (2**17)*0+(2**8)*111+115, (2**17)*0+(2**8)*112+168, (2**17)*0+(2**8)*165+  0, (2**17)*1+(2**8)*170+  4, 
(2**17)*0+(2**8)* 26+105, (2**17)*0+(2**8)* 26+ 70, (2**17)*0+(2**8)*111+151, (2**17)*0+(2**8)*125+ 29, (2**17)*0+(2**8)*129+115, (2**17)*0+(2**8)*137+132, (2**17)*0+(2**8)*157+  5, (2**17)*0+(2**8)*166+  0, (2**17)*1+(2**8)*210+118, 
(2**17)*0+(2**8)*  9+142, (2**17)*0+(2**8)* 19+144, (2**17)*0+(2**8)* 27+ 28, (2**17)*0+(2**8)* 27+ 38, (2**17)*0+(2**8)*109+118, (2**17)*0+(2**8)*135+ 55, (2**17)*0+(2**8)*150+133, (2**17)*0+(2**8)*167+  0, (2**17)*1+(2**8)*187+152, 
(2**17)*0+(2**8)* 62+138, (2**17)*0+(2**8)*109+178, (2**17)*0+(2**8)*114+ 62, (2**17)*0+(2**8)*128+ 31, (2**17)*0+(2**8)*129+169, (2**17)*0+(2**8)*138+153, (2**17)*0+(2**8)*143+ 17, (2**17)*0+(2**8)*168+  0, (2**17)*1+(2**8)*194+ 45, 
(2**17)*0+(2**8)* 17+103, (2**17)*0+(2**8)* 25+ 24, (2**17)*0+(2**8)* 76+157, (2**17)*0+(2**8)*109+139, (2**17)*0+(2**8)*109+120, (2**17)*0+(2**8)*119+ 88, (2**17)*0+(2**8)*140+142, (2**17)*0+(2**8)*159+ 92, (2**17)*1+(2**8)*169+  0, 
(2**17)*0+(2**8)*  0+ 21, (2**17)*0+(2**8)* 14+137, (2**17)*0+(2**8)* 35+ 10, (2**17)*0+(2**8)* 52+146, (2**17)*0+(2**8)*124+ 24, (2**17)*0+(2**8)*125+106, (2**17)*0+(2**8)*136+142, (2**17)*0+(2**8)*170+  0, (2**17)*1+(2**8)*184+ 48, 
(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  6+ 90, (2**17)*0+(2**8)* 10+103, (2**17)*0+(2**8)* 16+ 90, (2**17)*0+(2**8)* 32+ 25, (2**17)*0+(2**8)* 83+105, (2**17)*0+(2**8)*143+ 25, (2**17)*0+(2**8)*151+ 76, (2**17)*1+(2**8)*171+  0, 
(2**17)*0+(2**8)* 10+ 85, (2**17)*0+(2**8)* 18+ 66, (2**17)*0+(2**8)* 32+126, (2**17)*0+(2**8)* 47+ 50, (2**17)*0+(2**8)* 72+173, (2**17)*0+(2**8)*110+ 38, (2**17)*0+(2**8)*118+ 32, (2**17)*0+(2**8)*138+157, (2**17)*1+(2**8)*172+  0, 
(2**17)*0+(2**8)*  2+158, (2**17)*0+(2**8)* 11+155, (2**17)*0+(2**8)* 59+ 74, (2**17)*0+(2**8)*113+140, (2**17)*0+(2**8)*118+114, (2**17)*0+(2**8)*135+ 47, (2**17)*0+(2**8)*138+114, (2**17)*0+(2**8)*173+  0, (2**17)*1+(2**8)*183+147, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)*  8+120, (2**17)*0+(2**8)*  8+ 36, (2**17)*0+(2**8)* 13+101, (2**17)*0+(2**8)* 22+176, (2**17)*0+(2**8)* 29+164, (2**17)*0+(2**8)* 99+ 25, (2**17)*0+(2**8)*161+158, (2**17)*1+(2**8)*174+  0, 
(2**17)*0+(2**8)* 26+139, (2**17)*0+(2**8)* 32+ 37, (2**17)*0+(2**8)* 85+ 99, (2**17)*0+(2**8)*109+174, (2**17)*0+(2**8)*112+ 77, (2**17)*0+(2**8)*118+ 64, (2**17)*0+(2**8)*141+ 75, (2**17)*0+(2**8)*160+ 42, (2**17)*1+(2**8)*175+  0, 
(2**17)*0+(2**8)*  7+ 98, (2**17)*0+(2**8)* 21+  9, (2**17)*0+(2**8)* 22+ 67, (2**17)*0+(2**8)* 32+111, (2**17)*0+(2**8)*114+145, (2**17)*0+(2**8)*131+ 71, (2**17)*0+(2**8)*174+ 94, (2**17)*0+(2**8)*176+  0, (2**17)*1+(2**8)*196+ 61, 
(2**17)*0+(2**8)*  2+ 76, (2**17)*0+(2**8)*  3+163, (2**17)*0+(2**8)*  8+ 96, (2**17)*0+(2**8)* 14+166, (2**17)*0+(2**8)* 16+170, (2**17)*0+(2**8)* 30+167, (2**17)*0+(2**8)* 38+ 74, (2**17)*0+(2**8)*177+  0, (2**17)*1+(2**8)*191+ 78, 
(2**17)*0+(2**8)*  0+ 80, (2**17)*0+(2**8)* 43+131, (2**17)*0+(2**8)*100+ 57, (2**17)*0+(2**8)*111+ 36, (2**17)*0+(2**8)*114+ 47, (2**17)*0+(2**8)*127+ 92, (2**17)*0+(2**8)*131+119, (2**17)*0+(2**8)*131+ 41, (2**17)*1+(2**8)*178+  0, 
(2**17)*0+(2**8)* 24+165, (2**17)*0+(2**8)* 36+128, (2**17)*0+(2**8)* 96+120, (2**17)*0+(2**8)*108+  1, (2**17)*0+(2**8)*111+ 87, (2**17)*0+(2**8)*111+ 80, (2**17)*0+(2**8)*121+ 82, (2**17)*0+(2**8)*135+162, (2**17)*1+(2**8)*179+  0, 
(2**17)*0+(2**8)*  1+  5, (2**17)*0+(2**8)*  4+  7, (2**17)*0+(2**8)* 24+ 20, (2**17)*0+(2**8)* 26+146, (2**17)*0+(2**8)* 47+153, (2**17)*0+(2**8)*106+ 24, (2**17)*0+(2**8)*113+ 45, (2**17)*0+(2**8)*121+  5, (2**17)*1+(2**8)*180+  0, 
(2**17)*0+(2**8)*  1+ 80, (2**17)*0+(2**8)* 16+ 51, (2**17)*0+(2**8)* 17+167, (2**17)*0+(2**8)* 19+119, (2**17)*0+(2**8)* 24+ 50, (2**17)*0+(2**8)* 65+ 29, (2**17)*0+(2**8)*103+137, (2**17)*0+(2**8)*113+104, (2**17)*1+(2**8)*181+  0, 
(2**17)*0+(2**8)*  9+159, (2**17)*0+(2**8)* 11+126, (2**17)*0+(2**8)* 12+138, (2**17)*0+(2**8)* 44+138, (2**17)*0+(2**8)*133+162, (2**17)*0+(2**8)*142+133, (2**17)*0+(2**8)*143+ 96, (2**17)*0+(2**8)*182+  0, (2**17)*1+(2**8)*182+ 34, 
(2**17)*0+(2**8)* 15+ 51, (2**17)*0+(2**8)* 20+151, (2**17)*0+(2**8)* 22+ 59, (2**17)*0+(2**8)* 29+ 61, (2**17)*0+(2**8)* 30+ 27, (2**17)*0+(2**8)* 86+ 16, (2**17)*0+(2**8)*128+114, (2**17)*0+(2**8)*150+144, (2**17)*1+(2**8)*183+  0, 
(2**17)*0+(2**8)* 11+ 53, (2**17)*0+(2**8)* 15+  7, (2**17)*0+(2**8)* 20+106, (2**17)*0+(2**8)* 25+ 10, (2**17)*0+(2**8)*128+177, (2**17)*0+(2**8)*134+ 49, (2**17)*0+(2**8)*166+151, (2**17)*0+(2**8)*184+  0, (2**17)*1+(2**8)*212+ 84, 
(2**17)*0+(2**8)*  4+114, (2**17)*0+(2**8)* 25+133, (2**17)*0+(2**8)* 25+170, (2**17)*0+(2**8)* 93+ 93, (2**17)*0+(2**8)*117+ 20, (2**17)*0+(2**8)*138+ 36, (2**17)*0+(2**8)*142+173, (2**17)*0+(2**8)*157+ 77, (2**17)*1+(2**8)*185+  0, 
(2**17)*0+(2**8)*  2+ 78, (2**17)*0+(2**8)* 22+163, (2**17)*0+(2**8)* 40+ 92, (2**17)*0+(2**8)* 81+168, (2**17)*0+(2**8)*108+ 20, (2**17)*0+(2**8)*118+ 12, (2**17)*0+(2**8)*137+ 69, (2**17)*0+(2**8)*139+144, (2**17)*1+(2**8)*186+  0, 
(2**17)*0+(2**8)* 24+ 90, (2**17)*0+(2**8)*112+ 98, (2**17)*0+(2**8)*120+  8, (2**17)*0+(2**8)*126+ 56, (2**17)*0+(2**8)*142+ 78, (2**17)*0+(2**8)*142+ 16, (2**17)*0+(2**8)*177+136, (2**17)*0+(2**8)*187+  0, (2**17)*1+(2**8)*196+100, 
(2**17)*0+(2**8)*  8+ 27, (2**17)*0+(2**8)* 12+ 86, (2**17)*0+(2**8)* 20+ 99, (2**17)*0+(2**8)* 26+136, (2**17)*0+(2**8)*116+149, (2**17)*0+(2**8)*123+175, (2**17)*0+(2**8)*172+ 66, (2**17)*0+(2**8)*188+  0, (2**17)*1+(2**8)*190+ 97, 
(2**17)*0+(2**8)* 18+171, (2**17)*0+(2**8)* 30+ 53, (2**17)*0+(2**8)* 30+155, (2**17)*0+(2**8)* 55+134, (2**17)*0+(2**8)*110+ 21, (2**17)*0+(2**8)*117+ 39, (2**17)*0+(2**8)*141+ 59, (2**17)*0+(2**8)*189+  0, (2**17)*1+(2**8)*214+ 20, 
(2**17)*0+(2**8)* 33+ 44, (2**17)*0+(2**8)* 34+ 49, (2**17)*0+(2**8)* 65+121, (2**17)*0+(2**8)*116+172, (2**17)*0+(2**8)*116+ 15, (2**17)*0+(2**8)*132+ 91, (2**17)*0+(2**8)*132+166, (2**17)*0+(2**8)*185+ 52, (2**17)*1+(2**8)*190+  0, 
(2**17)*0+(2**8)*  7+ 62, (2**17)*0+(2**8)* 26+130, (2**17)*0+(2**8)* 35+ 19, (2**17)*0+(2**8)*121+ 25, (2**17)*0+(2**8)*129+162, (2**17)*0+(2**8)*134+ 39, (2**17)*0+(2**8)*162+137, (2**17)*0+(2**8)*191+  0, (2**17)*1+(2**8)*199+ 28, 
(2**17)*0+(2**8)*  4+145, (2**17)*0+(2**8)* 21+ 89, (2**17)*0+(2**8)* 72+ 96, (2**17)*0+(2**8)*120+131, (2**17)*0+(2**8)*121+159, (2**17)*0+(2**8)*129+177, (2**17)*0+(2**8)*135+155, (2**17)*0+(2**8)*179+120, (2**17)*1+(2**8)*192+  0, 
(2**17)*0+(2**8)* 13+ 89, (2**17)*0+(2**8)* 23+123, (2**17)*0+(2**8)*111+154, (2**17)*0+(2**8)*117+137, (2**17)*0+(2**8)*128+ 12, (2**17)*0+(2**8)*136+ 28, (2**17)*0+(2**8)*164+ 25, (2**17)*0+(2**8)*181+156, (2**17)*1+(2**8)*193+  0, 
(2**17)*0+(2**8)*  5+ 65, (2**17)*0+(2**8)*  7+116, (2**17)*0+(2**8)* 14+  5, (2**17)*0+(2**8)* 29+163, (2**17)*0+(2**8)* 32+ 68, (2**17)*0+(2**8)* 37+ 20, (2**17)*0+(2**8)*107+ 23, (2**17)*0+(2**8)*128+126, (2**17)*1+(2**8)*194+  0, 
(2**17)*0+(2**8)* 14+ 34, (2**17)*0+(2**8)* 23+ 37, (2**17)*0+(2**8)* 57+ 92, (2**17)*0+(2**8)* 84+107, (2**17)*0+(2**8)*109+156, (2**17)*0+(2**8)*120+139, (2**17)*0+(2**8)*141+132, (2**17)*0+(2**8)*142+172, (2**17)*1+(2**8)*195+  0, 
(2**17)*0+(2**8)* 21+ 58, (2**17)*0+(2**8)* 23+111, (2**17)*0+(2**8)* 33+ 72, (2**17)*0+(2**8)*115+ 38, (2**17)*0+(2**8)*122+ 61, (2**17)*0+(2**8)*129+ 28, (2**17)*0+(2**8)*147+ 54, (2**17)*0+(2**8)*195+173, (2**17)*1+(2**8)*196+  0, 
(2**17)*0+(2**8)*  0+138, (2**17)*0+(2**8)*  9+ 16, (2**17)*0+(2**8)* 61+ 25, (2**17)*0+(2**8)* 78+ 88, (2**17)*0+(2**8)*115+165, (2**17)*0+(2**8)*117+156, (2**17)*0+(2**8)*121+ 57, (2**17)*0+(2**8)*136+ 34, (2**17)*1+(2**8)*197+  0, 
(2**17)*0+(2**8)* 16+114, (2**17)*0+(2**8)* 16+101, (2**17)*0+(2**8)* 17+ 25, (2**17)*0+(2**8)* 19+175, (2**17)*0+(2**8)* 32+ 17, (2**17)*0+(2**8)*105+ 53, (2**17)*0+(2**8)*124+ 64, (2**17)*0+(2**8)*176+161, (2**17)*1+(2**8)*198+  0, 
(2**17)*0+(2**8)*  1+ 44, (2**17)*0+(2**8)* 12+145, (2**17)*0+(2**8)* 27+ 55, (2**17)*0+(2**8)* 29+ 91, (2**17)*0+(2**8)* 63+ 39, (2**17)*0+(2**8)*126+115, (2**17)*0+(2**8)*139+ 82, (2**17)*0+(2**8)*199+  0, (2**17)*1+(2**8)*209+139, 
(2**17)*0+(2**8)* 15+ 32, (2**17)*0+(2**8)* 18+172, (2**17)*0+(2**8)* 18+179, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 22+ 12, (2**17)*0+(2**8)* 68+ 80, (2**17)*0+(2**8)*124+ 25, (2**17)*0+(2**8)*200+  0, (2**17)*1+(2**8)*213+158, 
(2**17)*0+(2**8)*  2+119, (2**17)*0+(2**8)* 12+ 42, (2**17)*0+(2**8)* 16+109, (2**17)*0+(2**8)* 19+ 25, (2**17)*0+(2**8)*117+132, (2**17)*0+(2**8)*142+ 50, (2**17)*0+(2**8)*169+ 44, (2**17)*0+(2**8)*193+ 65, (2**17)*1+(2**8)*201+  0, 
(2**17)*0+(2**8)* 95+ 10, (2**17)*0+(2**8)*108+ 71, (2**17)*0+(2**8)*113+  7, (2**17)*0+(2**8)*133+122, (2**17)*0+(2**8)*136+ 50, (2**17)*0+(2**8)*139+ 55, (2**17)*0+(2**8)*142+ 20, (2**17)*0+(2**8)*175+ 12, (2**17)*1+(2**8)*202+  0, 
(2**17)*0+(2**8)*  5+ 98, (2**17)*0+(2**8)* 16+164, (2**17)*0+(2**8)*111+176, (2**17)*0+(2**8)*112+ 74, (2**17)*0+(2**8)*120+166, (2**17)*0+(2**8)*127+ 35, (2**17)*0+(2**8)*147+ 85, (2**17)*0+(2**8)*182+ 87, (2**17)*1+(2**8)*203+  0, 
(2**17)*0+(2**8)*  2+ 99, (2**17)*0+(2**8)* 28+ 48, (2**17)*0+(2**8)* 80+  7, (2**17)*0+(2**8)*114+154, (2**17)*0+(2**8)*133+125, (2**17)*0+(2**8)*141+ 79, (2**17)*0+(2**8)*143+104, (2**17)*0+(2**8)*179+ 95, (2**17)*1+(2**8)*204+  0, 
(2**17)*0+(2**8)*  3+136, (2**17)*0+(2**8)*  5+115, (2**17)*0+(2**8)* 14+168, (2**17)*0+(2**8)* 20+ 86, (2**17)*0+(2**8)* 21+154, (2**17)*0+(2**8)* 50+ 95, (2**17)*0+(2**8)*126+141, (2**17)*0+(2**8)*205+  0, (2**17)*1+(2**8)*208+  9, 
(2**17)*0+(2**8)* 33+113, (2**17)*0+(2**8)* 37+ 72, (2**17)*0+(2**8)*108+ 57, (2**17)*0+(2**8)*120+ 30, (2**17)*0+(2**8)*137+148, (2**17)*0+(2**8)*138+ 92, (2**17)*0+(2**8)*140+ 78, (2**17)*0+(2**8)*192+ 32, (2**17)*1+(2**8)*206+  0, 
(2**17)*0+(2**8)*  1+156, (2**17)*0+(2**8)* 28+169, (2**17)*0+(2**8)* 31+178, (2**17)*0+(2**8)* 66+156, (2**17)*0+(2**8)*112+ 39, (2**17)*0+(2**8)*130+174, (2**17)*0+(2**8)*140+158, (2**17)*0+(2**8)*181+ 46, (2**17)*1+(2**8)*207+  0, 
(2**17)*0+(2**8)*  6+ 47, (2**17)*0+(2**8)*  8+114, (2**17)*0+(2**8)* 23+146, (2**17)*0+(2**8)* 34+112, (2**17)*0+(2**8)* 35+160, (2**17)*0+(2**8)*118+ 76, (2**17)*0+(2**8)*153+ 78, (2**17)*0+(2**8)*186+169, (2**17)*1+(2**8)*208+  0, 
(2**17)*0+(2**8)*  7+136, (2**17)*0+(2**8)* 14+ 76, (2**17)*0+(2**8)* 17+117, (2**17)*0+(2**8)*107+ 53, (2**17)*0+(2**8)*134+ 97, (2**17)*0+(2**8)*139+118, (2**17)*0+(2**8)*143+ 41, (2**17)*0+(2**8)*178+ 94, (2**17)*1+(2**8)*209+  0, 
(2**17)*0+(2**8)*  5+  9, (2**17)*0+(2**8)* 19+170, (2**17)*0+(2**8)*128+121, (2**17)*0+(2**8)*129+ 44, (2**17)*0+(2**8)*132+170, (2**17)*0+(2**8)*137+ 98, (2**17)*0+(2**8)*178+ 93, (2**17)*0+(2**8)*195+171, (2**17)*1+(2**8)*210+  0, 
(2**17)*0+(2**8)*  6+108, (2**17)*0+(2**8)*  6+149, (2**17)*0+(2**8)* 10+ 18, (2**17)*0+(2**8)* 28+ 73, (2**17)*0+(2**8)* 33+ 39, (2**17)*0+(2**8)* 34+ 87, (2**17)*0+(2**8)* 89+  8, (2**17)*0+(2**8)*154+143, (2**17)*1+(2**8)*211+  0, 
(2**17)*0+(2**8)*  5+ 59, (2**17)*0+(2**8)* 14+ 55, (2**17)*0+(2**8)* 17+157, (2**17)*0+(2**8)* 26+ 86, (2**17)*0+(2**8)* 95+ 41, (2**17)*0+(2**8)*112+108, (2**17)*0+(2**8)*114+  3, (2**17)*0+(2**8)*161+ 40, (2**17)*1+(2**8)*212+  0, 
(2**17)*0+(2**8)* 11+176, (2**17)*0+(2**8)* 35+  3, (2**17)*0+(2**8)* 48+152, (2**17)*0+(2**8)*120+172, (2**17)*0+(2**8)*126+ 93, (2**17)*0+(2**8)*127+142, (2**17)*0+(2**8)*136+ 99, (2**17)*0+(2**8)*201+ 42, (2**17)*1+(2**8)*213+  0, 
(2**17)*0+(2**8)* 16+155, (2**17)*0+(2**8)* 28+ 29, (2**17)*0+(2**8)*121+ 77, (2**17)*0+(2**8)*127+ 68, (2**17)*0+(2**8)*132+137, (2**17)*0+(2**8)*136+  7, (2**17)*0+(2**8)*154+104, (2**17)*0+(2**8)*198+144, (2**17)*1+(2**8)*214+  0, 
(2**17)*0+(2**8)* 21+144, (2**17)*0+(2**8)* 31+170, (2**17)*0+(2**8)* 98+142, (2**17)*0+(2**8)*118+  5, (2**17)*0+(2**8)*123+ 38, (2**17)*0+(2**8)*127+ 98, (2**17)*0+(2**8)*129+ 56, (2**17)*0+(2**8)*162+ 29, (2**17)*1+(2**8)*215+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  0+  2, (2**17)*0+(2**8)* 11+118, (2**17)*0+(2**8)* 12+115, (2**17)*0+(2**8)* 39+142, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 79+116, (2**17)*1+(2**8)*199+ 83, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 12+118, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)*112+151, (2**17)*0+(2**8)*123+ 95, (2**17)*0+(2**8)*127+156, (2**17)*0+(2**8)*137+113, (2**17)*1+(2**8)*231+ 31, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 11+ 36, (2**17)*0+(2**8)* 39+159, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 85+ 36, (2**17)*0+(2**8)*117+ 56, (2**17)*0+(2**8)*128+ 76, (2**17)*1+(2**8)*167+176, 
(2**17)*0+(2**8)*  1+154, (2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)*114+150, (2**17)*0+(2**8)*123+ 52, (2**17)*0+(2**8)*126+115, (2**17)*0+(2**8)*136+ 10, (2**17)*1+(2**8)*226+134, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 72+133, (2**17)*0+(2**8)* 78+ 17, (2**17)*0+(2**8)*121+ 49, (2**17)*0+(2**8)*122+101, (2**17)*0+(2**8)*150+170, (2**17)*1+(2**8)*178+ 16, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  5+156, (2**17)*0+(2**8)*  7+ 46, (2**17)*0+(2**8)*  9+ 79, (2**17)*0+(2**8)* 57+ 82, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)*182+ 26, (2**17)*1+(2**8)*186+ 97, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  6+  4, (2**17)*0+(2**8)* 35+ 48, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 69+ 10, (2**17)*0+(2**8)* 83+ 81, (2**17)*0+(2**8)*120+ 69, (2**17)*1+(2**8)*128+107, 
(2**17)*0+(2**8)*  0+ 23, (2**17)*0+(2**8)*  1+112, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  7+172, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 99+143, (2**17)*0+(2**8)*134+134, (2**17)*1+(2**8)*208+ 62, 
(2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 10+  3, (2**17)*0+(2**8)* 11+105, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)*107+ 42, (2**17)*0+(2**8)*133+ 25, (2**17)*0+(2**8)*151+122, (2**17)*1+(2**8)*230+135, 
(2**17)*0+(2**8)*  4+164, (2**17)*0+(2**8)*  5+103, (2**17)*0+(2**8)*  7+ 88, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 42+ 52, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 94+ 13, (2**17)*1+(2**8)*223+154, 
(2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 38+ 34, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)*126+104, (2**17)*0+(2**8)*127+ 68, (2**17)*0+(2**8)*162+159, (2**17)*0+(2**8)*205+ 67, (2**17)*1+(2**8)*214+ 63, 
(2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 33+162, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 82+ 51, (2**17)*0+(2**8)*122+ 60, (2**17)*0+(2**8)*126+ 47, (2**17)*0+(2**8)*128+ 32, (2**17)*1+(2**8)*217+  2, 
(2**17)*0+(2**8)*  3+ 83, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 44+ 98, (2**17)*0+(2**8)* 56+ 20, (2**17)*0+(2**8)* 63+152, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)*129+169, (2**17)*1+(2**8)*223+ 71, 
(2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)* 76+  2, (2**17)*0+(2**8)*120+156, (2**17)*0+(2**8)*121+ 54, (2**17)*0+(2**8)*131+ 34, (2**17)*0+(2**8)*160+169, (2**17)*1+(2**8)*185+ 85, 
(2**17)*0+(2**8)*  4+149, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 23+105, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 82+ 45, (2**17)*0+(2**8)*122+107, (2**17)*0+(2**8)*147+137, (2**17)*1+(2**8)*197+ 11, 
(2**17)*0+(2**8)*  2+ 37, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 56+144, (2**17)*0+(2**8)* 71+ 78, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)*130+  8, (2**17)*0+(2**8)*145+147, (2**17)*1+(2**8)*227+147, 
(2**17)*0+(2**8)*  3+121, (2**17)*0+(2**8)* 10+113, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 34+  4, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)* 86+130, (2**17)*0+(2**8)*102+ 42, (2**17)*1+(2**8)*139+180, 
(2**17)*0+(2**8)*  6+ 96, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 34+ 35, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)* 78+123, (2**17)*0+(2**8)*108+ 40, (2**17)*0+(2**8)*122+150, (2**17)*1+(2**8)*125+ 17, 
(2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)*125+127, (2**17)*0+(2**8)*129+138, (2**17)*0+(2**8)*149+ 56, (2**17)*0+(2**8)*158+ 49, (2**17)*0+(2**8)*186+ 76, (2**17)*1+(2**8)*208+173, 
(2**17)*0+(2**8)*  0+ 88, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 47+ 98, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)*129+167, (2**17)*0+(2**8)*170+ 28, (2**17)*0+(2**8)*187+ 45, (2**17)*1+(2**8)*204+ 46, 
(2**17)*0+(2**8)*  5+ 14, (2**17)*0+(2**8)* 16+ 75, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 61+ 78, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)*121+ 43, (2**17)*0+(2**8)*164+165, (2**17)*1+(2**8)*210+ 22, 
(2**17)*0+(2**8)*  7+101, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 28+ 58, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)*127+154, (2**17)*0+(2**8)*156+ 88, (2**17)*0+(2**8)*201+ 83, (2**17)*1+(2**8)*207+130, 
(2**17)*0+(2**8)*  3+ 68, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 55+ 43, (2**17)*0+(2**8)* 70+  9, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)*128+ 81, (2**17)*0+(2**8)*168+ 81, (2**17)*1+(2**8)*194+ 67, 
(2**17)*0+(2**8)*  4+ 51, (2**17)*0+(2**8)* 11+ 85, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)*115+ 44, (2**17)*0+(2**8)*120+134, (2**17)*0+(2**8)*173+ 50, (2**17)*1+(2**8)*235+ 26, 
(2**17)*0+(2**8)*  2+ 50, (2**17)*0+(2**8)*  8+127, (2**17)*0+(2**8)* 11+179, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 68+ 75, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)*165+164, (2**17)*1+(2**8)*209+157, 
(2**17)*0+(2**8)*  0+ 67, (2**17)*0+(2**8)*  1+115, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 37+ 99, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*105+136, (2**17)*0+(2**8)*129+163, (2**17)*1+(2**8)*218+156, 
(2**17)*0+(2**8)*  0+  4, (2**17)*0+(2**8)*  4+ 44, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 54+ 61, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)*174+ 98, (2**17)*0+(2**8)*197+161, (2**17)*1+(2**8)*201+152, 
(2**17)*0+(2**8)*  1+143, (2**17)*0+(2**8)*  4+139, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 30+108, (2**17)*0+(2**8)* 72+ 50, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)* 96+ 76, (2**17)*1+(2**8)*178+ 56, 
(2**17)*0+(2**8)*  2+155, (2**17)*0+(2**8)* 10+ 38, (2**17)*0+(2**8)* 10+ 29, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)*105+106, (2**17)*0+(2**8)*142+ 84, (2**17)*1+(2**8)*233+ 75, 
(2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 73+123, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)* 91+149, (2**17)*0+(2**8)*129+ 77, (2**17)*0+(2**8)*131+ 69, (2**17)*0+(2**8)*148+ 62, (2**17)*1+(2**8)*175+ 47, 
(2**17)*0+(2**8)* 18+ 18, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 86+ 46, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)*125+141, (2**17)*0+(2**8)*129+ 56, (2**17)*0+(2**8)*155+ 61, (2**17)*1+(2**8)*217+139, 
(2**17)*0+(2**8)*  6+145, (2**17)*0+(2**8)*  7+119, (2**17)*0+(2**8)* 11+  5, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)*100+ 28, (2**17)*0+(2**8)*124+ 39, (2**17)*1+(2**8)*237+ 40, 
(2**17)*0+(2**8)*  5+ 21, (2**17)*0+(2**8)*  7+ 68, (2**17)*0+(2**8)* 11+117, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*121+107, (2**17)*0+(2**8)*193+ 54, (2**17)*1+(2**8)*200+  4, 
(2**17)*0+(2**8)*  1+ 69, (2**17)*0+(2**8)*  9+ 61, (2**17)*0+(2**8)* 10+ 92, (2**17)*0+(2**8)* 26+ 49, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*113+ 98, (2**17)*1+(2**8)*224+101, 
(2**17)*0+(2**8)*  3+145, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 65+ 89, (2**17)*0+(2**8)* 69+136, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*127+ 98, (2**17)*0+(2**8)*172+ 66, (2**17)*1+(2**8)*177+171, 
(2**17)*0+(2**8)*  2+ 49, (2**17)*0+(2**8)* 11+103, (2**17)*0+(2**8)* 23+  4, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 68+ 79, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*108+158, (2**17)*1+(2**8)*146+ 71, 
(2**17)*0+(2**8)*  3+ 46, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 51+ 36, (2**17)*0+(2**8)* 71+173, (2**17)*0+(2**8)* 91+ 54, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*125+101, (2**17)*1+(2**8)*139+102, 
(2**17)*0+(2**8)*  2+170, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)* 99+174, (2**17)*0+(2**8)*123+165, (2**17)*0+(2**8)*129+ 65, (2**17)*0+(2**8)*140+166, (2**17)*1+(2**8)*218+130, 
(2**17)*0+(2**8)* 21+ 66, (2**17)*0+(2**8)* 32+149, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*124+122, (2**17)*0+(2**8)*129+ 70, (2**17)*0+(2**8)*212+  1, (2**17)*1+(2**8)*222+ 77, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*0+(2**8)* 11+166, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 93+171, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*111+ 25, (2**17)*0+(2**8)*149+133, (2**17)*1+(2**8)*157+170, 
(2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 53+ 36, (2**17)*0+(2**8)* 95+133, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*118+ 66, (2**17)*0+(2**8)*121+ 83, (2**17)*0+(2**8)*127+ 35, (2**17)*1+(2**8)*142+133, 
(2**17)*0+(2**8)*  2+ 72, (2**17)*0+(2**8)*  7+131, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 46+ 29, (2**17)*0+(2**8)* 64+ 76, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*144+ 71, (2**17)*1+(2**8)*207+ 89, 
(2**17)*0+(2**8)*  5+132, (2**17)*0+(2**8)* 10+168, (2**17)*0+(2**8)* 15+ 92, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 64+130, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*168+109, (2**17)*1+(2**8)*195+123, 
(2**17)*0+(2**8)*  6+ 12, (2**17)*0+(2**8)*  9+ 26, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*109+137, (2**17)*0+(2**8)*147+ 87, (2**17)*0+(2**8)*153+ 56, (2**17)*1+(2**8)*216+ 86, 
(2**17)*0+(2**8)*  4+172, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 59+171, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*121+ 52, (2**17)*0+(2**8)*145+140, (2**17)*0+(2**8)*210+ 75, (2**17)*1+(2**8)*213+ 31, 
(2**17)*0+(2**8)* 36+ 74, (2**17)*0+(2**8)* 41+161, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 76+ 25, (2**17)*0+(2**8)* 84+100, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*126+118, (2**17)*1+(2**8)*130+ 91, 
(2**17)*0+(2**8)*  8+160, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*120+107, (2**17)*0+(2**8)*135+171, (2**17)*0+(2**8)*161+163, (2**17)*0+(2**8)*180+152, (2**17)*1+(2**8)*181+ 69, 
(2**17)*0+(2**8)*  6+ 32, (2**17)*0+(2**8)* 13+ 80, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 50+ 92, (2**17)*0+(2**8)* 60+143, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*126+127, (2**17)*1+(2**8)*234+112, 
(2**17)*0+(2**8)*  0+174, (2**17)*0+(2**8)*  4+ 13, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*138+ 13, (2**17)*0+(2**8)*165+ 62, (2**17)*0+(2**8)*212+ 93, (2**17)*1+(2**8)*236+139, 
(2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 75+117, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*123+148, (2**17)*0+(2**8)*125+ 26, (2**17)*0+(2**8)*130+ 56, (2**17)*0+(2**8)*141+ 35, (2**17)*1+(2**8)*239+ 30, 
(2**17)*0+(2**8)*  2+ 91, (2**17)*0+(2**8)*  8+ 83, (2**17)*0+(2**8)* 24+ 70, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*112+158, (2**17)*0+(2**8)*151+ 21, (2**17)*1+(2**8)*239+122, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*0+(2**8)*  5+ 40, (2**17)*0+(2**8)* 10+176, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*116+  4, (2**17)*0+(2**8)*126+ 51, (2**17)*1+(2**8)*194+155, 
(2**17)*0+(2**8)*  3+154, (2**17)*0+(2**8)*  8+ 84, (2**17)*0+(2**8)* 51+157, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 95+ 97, (2**17)*0+(2**8)*101+167, (2**17)*0+(2**8)*112+  0, (2**17)*1+(2**8)*160+103, 
(2**17)*0+(2**8)* 14+122, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*126+ 62, (2**17)*0+(2**8)*130+137, (2**17)*0+(2**8)*163+160, (2**17)*0+(2**8)*182+ 59, (2**17)*1+(2**8)*224+173, 
(2**17)*0+(2**8)*  8+ 45, (2**17)*0+(2**8)* 11+162, (2**17)*0+(2**8)* 17+ 33, (2**17)*0+(2**8)* 49+ 74, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 80+ 61, (2**17)*0+(2**8)*114+  0, (2**17)*1+(2**8)*190+125, 
(2**17)*0+(2**8)*  4+119, (2**17)*0+(2**8)* 20+ 17, (2**17)*0+(2**8)* 32+ 55, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)*106+ 92, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*118+ 47, (2**17)*1+(2**8)*128+ 89, 
(2**17)*0+(2**8)*  2+121, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 59+ 43, (2**17)*0+(2**8)*100+ 35, (2**17)*0+(2**8)*109+ 29, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*129+  6, (2**17)*1+(2**8)*166+134, 
(2**17)*0+(2**8)* 49+ 43, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*123+129, (2**17)*0+(2**8)*130+ 36, (2**17)*0+(2**8)*163+ 92, (2**17)*0+(2**8)*183+112, (2**17)*1+(2**8)*203+ 84, 
(2**17)*0+(2**8)*  4+ 25, (2**17)*0+(2**8)*  5+ 81, (2**17)*0+(2**8)* 52+ 32, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 67+ 78, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*128+166, (2**17)*1+(2**8)*209+ 21, 
(2**17)*0+(2**8)*  1+148, (2**17)*0+(2**8)*  3+ 36, (2**17)*0+(2**8)*  4+  5, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)*101+143, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*128+123, (2**17)*1+(2**8)*230+ 12, 
(2**17)*0+(2**8)* 79+ 82, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*120+  2, (2**17)*0+(2**8)*131+118, (2**17)*0+(2**8)*132+115, (2**17)*0+(2**8)*159+142, (2**17)*0+(2**8)*180+  0, (2**17)*1+(2**8)*199+116, 
(2**17)*0+(2**8)*  3+ 94, (2**17)*0+(2**8)*  7+155, (2**17)*0+(2**8)* 17+112, (2**17)*0+(2**8)*111+ 30, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*132+118, (2**17)*0+(2**8)*181+  0, (2**17)*1+(2**8)*232+151, 
(2**17)*0+(2**8)*  8+ 75, (2**17)*0+(2**8)* 47+175, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*131+ 36, (2**17)*0+(2**8)*159+159, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*205+ 36, (2**17)*1+(2**8)*237+ 56, 
(2**17)*0+(2**8)*  3+ 51, (2**17)*0+(2**8)*  6+114, (2**17)*0+(2**8)* 16+  9, (2**17)*0+(2**8)*106+133, (2**17)*0+(2**8)*121+154, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*183+  0, (2**17)*1+(2**8)*234+150, 
(2**17)*0+(2**8)*  1+ 48, (2**17)*0+(2**8)*  2+100, (2**17)*0+(2**8)* 30+169, (2**17)*0+(2**8)* 58+ 15, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*192+133, (2**17)*1+(2**8)*198+ 17, 
(2**17)*0+(2**8)* 62+ 25, (2**17)*0+(2**8)* 66+ 96, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*125+156, (2**17)*0+(2**8)*127+ 46, (2**17)*0+(2**8)*129+ 79, (2**17)*0+(2**8)*177+ 82, (2**17)*1+(2**8)*185+  0, 
(2**17)*0+(2**8)*  0+ 68, (2**17)*0+(2**8)*  8+106, (2**17)*0+(2**8)*126+  0, (2**17)*0+(2**8)*126+  4, (2**17)*0+(2**8)*155+ 48, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*189+ 10, (2**17)*1+(2**8)*203+ 81, 
(2**17)*0+(2**8)* 14+133, (2**17)*0+(2**8)* 88+ 61, (2**17)*0+(2**8)*120+ 23, (2**17)*0+(2**8)*121+112, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*127+172, (2**17)*0+(2**8)*187+  0, (2**17)*1+(2**8)*219+143, 
(2**17)*0+(2**8)* 13+ 24, (2**17)*0+(2**8)* 31+121, (2**17)*0+(2**8)*110+134, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*130+  3, (2**17)*0+(2**8)*131+105, (2**17)*0+(2**8)*188+  0, (2**17)*1+(2**8)*227+ 42, 
(2**17)*0+(2**8)*103+153, (2**17)*0+(2**8)*124+164, (2**17)*0+(2**8)*125+103, (2**17)*0+(2**8)*127+ 88, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*162+ 52, (2**17)*0+(2**8)*189+  0, (2**17)*1+(2**8)*214+ 13, 
(2**17)*0+(2**8)*  6+103, (2**17)*0+(2**8)*  7+ 67, (2**17)*0+(2**8)* 42+158, (2**17)*0+(2**8)* 85+ 66, (2**17)*0+(2**8)* 94+ 62, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*158+ 34, (2**17)*1+(2**8)*190+  0, 
(2**17)*0+(2**8)*  2+ 59, (2**17)*0+(2**8)*  6+ 46, (2**17)*0+(2**8)*  8+ 31, (2**17)*0+(2**8)* 97+  1, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*153+162, (2**17)*0+(2**8)*191+  0, (2**17)*1+(2**8)*202+ 51, 
(2**17)*0+(2**8)*  9+168, (2**17)*0+(2**8)*103+ 70, (2**17)*0+(2**8)*123+ 83, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*164+ 98, (2**17)*0+(2**8)*176+ 20, (2**17)*0+(2**8)*183+152, (2**17)*1+(2**8)*192+  0, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)*  1+ 53, (2**17)*0+(2**8)* 11+ 33, (2**17)*0+(2**8)* 40+168, (2**17)*0+(2**8)* 65+ 84, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*193+  0, (2**17)*1+(2**8)*196+  2, 
(2**17)*0+(2**8)*  2+106, (2**17)*0+(2**8)* 27+136, (2**17)*0+(2**8)* 77+ 10, (2**17)*0+(2**8)*124+149, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*143+105, (2**17)*0+(2**8)*194+  0, (2**17)*1+(2**8)*202+ 45, 
(2**17)*0+(2**8)* 10+  7, (2**17)*0+(2**8)* 25+146, (2**17)*0+(2**8)*107+146, (2**17)*0+(2**8)*122+ 37, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*176+144, (2**17)*0+(2**8)*191+ 78, (2**17)*1+(2**8)*195+  0, 
(2**17)*0+(2**8)* 19+179, (2**17)*0+(2**8)*123+121, (2**17)*0+(2**8)*130+113, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*154+  4, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*206+130, (2**17)*1+(2**8)*222+ 42, 
(2**17)*0+(2**8)*  2+149, (2**17)*0+(2**8)*  5+ 16, (2**17)*0+(2**8)*126+ 96, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*154+ 35, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*198+123, (2**17)*1+(2**8)*228+ 40, 
(2**17)*0+(2**8)*  5+126, (2**17)*0+(2**8)*  9+137, (2**17)*0+(2**8)* 29+ 55, (2**17)*0+(2**8)* 38+ 48, (2**17)*0+(2**8)* 66+ 75, (2**17)*0+(2**8)* 88+172, (2**17)*0+(2**8)*138+  0, (2**17)*1+(2**8)*198+  0, 
(2**17)*0+(2**8)*  9+166, (2**17)*0+(2**8)* 50+ 27, (2**17)*0+(2**8)* 67+ 44, (2**17)*0+(2**8)* 84+ 45, (2**17)*0+(2**8)*120+ 88, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*167+ 98, (2**17)*1+(2**8)*199+  0, 
(2**17)*0+(2**8)*  1+ 42, (2**17)*0+(2**8)* 44+164, (2**17)*0+(2**8)* 90+ 21, (2**17)*0+(2**8)*125+ 14, (2**17)*0+(2**8)*136+ 75, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*181+ 78, (2**17)*1+(2**8)*200+  0, 
(2**17)*0+(2**8)*  7+153, (2**17)*0+(2**8)* 36+ 87, (2**17)*0+(2**8)* 81+ 82, (2**17)*0+(2**8)* 87+129, (2**17)*0+(2**8)*127+101, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*148+ 58, (2**17)*1+(2**8)*201+  0, 
(2**17)*0+(2**8)*  8+ 80, (2**17)*0+(2**8)* 48+ 80, (2**17)*0+(2**8)* 74+ 66, (2**17)*0+(2**8)*123+ 68, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*175+ 43, (2**17)*0+(2**8)*190+  9, (2**17)*1+(2**8)*202+  0, 
(2**17)*0+(2**8)*  0+133, (2**17)*0+(2**8)* 53+ 49, (2**17)*0+(2**8)*115+ 25, (2**17)*0+(2**8)*124+ 51, (2**17)*0+(2**8)*131+ 85, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*203+  0, (2**17)*1+(2**8)*235+ 44, 
(2**17)*0+(2**8)* 45+163, (2**17)*0+(2**8)* 89+156, (2**17)*0+(2**8)*122+ 50, (2**17)*0+(2**8)*128+127, (2**17)*0+(2**8)*131+179, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*188+ 75, (2**17)*1+(2**8)*204+  0, 
(2**17)*0+(2**8)*  9+162, (2**17)*0+(2**8)* 98+155, (2**17)*0+(2**8)*120+ 67, (2**17)*0+(2**8)*121+115, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*157+ 99, (2**17)*0+(2**8)*205+  0, (2**17)*1+(2**8)*225+136, 
(2**17)*0+(2**8)* 54+ 97, (2**17)*0+(2**8)* 77+160, (2**17)*0+(2**8)* 81+151, (2**17)*0+(2**8)*120+  4, (2**17)*0+(2**8)*124+ 44, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*174+ 61, (2**17)*1+(2**8)*206+  0, 
(2**17)*0+(2**8)* 58+ 55, (2**17)*0+(2**8)*121+143, (2**17)*0+(2**8)*124+139, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*150+108, (2**17)*0+(2**8)*192+ 50, (2**17)*0+(2**8)*207+  0, (2**17)*1+(2**8)*216+ 76, 
(2**17)*0+(2**8)* 22+ 83, (2**17)*0+(2**8)*113+ 74, (2**17)*0+(2**8)*122+155, (2**17)*0+(2**8)*130+ 38, (2**17)*0+(2**8)*130+ 29, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*208+  0, (2**17)*1+(2**8)*225+106, 
(2**17)*0+(2**8)*  9+ 76, (2**17)*0+(2**8)* 11+ 68, (2**17)*0+(2**8)* 28+ 61, (2**17)*0+(2**8)* 55+ 46, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*193+123, (2**17)*0+(2**8)*209+  0, (2**17)*1+(2**8)*211+149, 
(2**17)*0+(2**8)*  5+140, (2**17)*0+(2**8)*  9+ 55, (2**17)*0+(2**8)* 35+ 60, (2**17)*0+(2**8)* 97+138, (2**17)*0+(2**8)*138+ 18, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*206+ 46, (2**17)*1+(2**8)*210+  0, 
(2**17)*0+(2**8)*  4+ 38, (2**17)*0+(2**8)*117+ 39, (2**17)*0+(2**8)*126+145, (2**17)*0+(2**8)*127+119, (2**17)*0+(2**8)*131+  5, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*211+  0, (2**17)*1+(2**8)*220+ 28, 
(2**17)*0+(2**8)*  1+106, (2**17)*0+(2**8)* 73+ 53, (2**17)*0+(2**8)* 80+  3, (2**17)*0+(2**8)*125+ 21, (2**17)*0+(2**8)*127+ 68, (2**17)*0+(2**8)*131+117, (2**17)*0+(2**8)*152+  0, (2**17)*1+(2**8)*212+  0, 
(2**17)*0+(2**8)*104+100, (2**17)*0+(2**8)*121+ 69, (2**17)*0+(2**8)*129+ 61, (2**17)*0+(2**8)*130+ 92, (2**17)*0+(2**8)*146+ 49, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*213+  0, (2**17)*1+(2**8)*233+ 98, 
(2**17)*0+(2**8)*  7+ 97, (2**17)*0+(2**8)* 52+ 65, (2**17)*0+(2**8)* 57+170, (2**17)*0+(2**8)*123+145, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*185+ 89, (2**17)*0+(2**8)*189+136, (2**17)*1+(2**8)*214+  0, 
(2**17)*0+(2**8)* 26+ 70, (2**17)*0+(2**8)*122+ 49, (2**17)*0+(2**8)*131+103, (2**17)*0+(2**8)*143+  4, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*188+ 79, (2**17)*0+(2**8)*215+  0, (2**17)*1+(2**8)*228+158, 
(2**17)*0+(2**8)*  5+100, (2**17)*0+(2**8)* 19+101, (2**17)*0+(2**8)*123+ 46, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*171+ 36, (2**17)*0+(2**8)*191+173, (2**17)*0+(2**8)*211+ 54, (2**17)*1+(2**8)*216+  0, 
(2**17)*0+(2**8)*  3+164, (2**17)*0+(2**8)*  9+ 64, (2**17)*0+(2**8)* 20+165, (2**17)*0+(2**8)* 98+129, (2**17)*0+(2**8)*122+170, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*217+  0, (2**17)*1+(2**8)*219+174, 
(2**17)*0+(2**8)*  4+121, (2**17)*0+(2**8)*  9+ 69, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*102+ 76, (2**17)*0+(2**8)*141+ 66, (2**17)*0+(2**8)*152+149, (2**17)*0+(2**8)*158+  0, (2**17)*1+(2**8)*218+  0, 
(2**17)*0+(2**8)* 29+132, (2**17)*0+(2**8)* 37+169, (2**17)*0+(2**8)*120+ 77, (2**17)*0+(2**8)*131+166, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*213+171, (2**17)*0+(2**8)*219+  0, (2**17)*1+(2**8)*231+ 25, 
(2**17)*0+(2**8)*  1+ 82, (2**17)*0+(2**8)*  7+ 34, (2**17)*0+(2**8)* 22+132, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*173+ 36, (2**17)*0+(2**8)*215+133, (2**17)*0+(2**8)*220+  0, (2**17)*1+(2**8)*238+ 66, 
(2**17)*0+(2**8)* 24+ 70, (2**17)*0+(2**8)* 87+ 88, (2**17)*0+(2**8)*122+ 72, (2**17)*0+(2**8)*127+131, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*166+ 29, (2**17)*0+(2**8)*184+ 76, (2**17)*1+(2**8)*221+  0, 
(2**17)*0+(2**8)* 48+108, (2**17)*0+(2**8)* 75+122, (2**17)*0+(2**8)*125+132, (2**17)*0+(2**8)*130+168, (2**17)*0+(2**8)*135+ 92, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*184+130, (2**17)*1+(2**8)*222+  0, 
(2**17)*0+(2**8)* 27+ 86, (2**17)*0+(2**8)* 33+ 55, (2**17)*0+(2**8)* 96+ 85, (2**17)*0+(2**8)*126+ 12, (2**17)*0+(2**8)*129+ 26, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*223+  0, (2**17)*1+(2**8)*229+137, 
(2**17)*0+(2**8)*  1+ 51, (2**17)*0+(2**8)* 25+139, (2**17)*0+(2**8)* 90+ 74, (2**17)*0+(2**8)* 93+ 30, (2**17)*0+(2**8)*124+172, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*179+171, (2**17)*1+(2**8)*224+  0, 
(2**17)*0+(2**8)*  6+117, (2**17)*0+(2**8)* 10+ 90, (2**17)*0+(2**8)*156+ 74, (2**17)*0+(2**8)*161+161, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*196+ 25, (2**17)*0+(2**8)*204+100, (2**17)*1+(2**8)*225+  0, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)* 15+170, (2**17)*0+(2**8)* 41+162, (2**17)*0+(2**8)* 60+151, (2**17)*0+(2**8)* 61+ 68, (2**17)*0+(2**8)*128+160, (2**17)*0+(2**8)*166+  0, (2**17)*1+(2**8)*226+  0, 
(2**17)*0+(2**8)*  6+126, (2**17)*0+(2**8)*114+111, (2**17)*0+(2**8)*126+ 32, (2**17)*0+(2**8)*133+ 80, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*170+ 92, (2**17)*0+(2**8)*180+143, (2**17)*1+(2**8)*227+  0, 
(2**17)*0+(2**8)* 18+ 12, (2**17)*0+(2**8)* 45+ 61, (2**17)*0+(2**8)* 92+ 92, (2**17)*0+(2**8)*116+138, (2**17)*0+(2**8)*120+174, (2**17)*0+(2**8)*124+ 13, (2**17)*0+(2**8)*168+  0, (2**17)*1+(2**8)*228+  0, 
(2**17)*0+(2**8)*  3+147, (2**17)*0+(2**8)*  5+ 25, (2**17)*0+(2**8)* 10+ 55, (2**17)*0+(2**8)* 21+ 34, (2**17)*0+(2**8)*119+ 29, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*195+117, (2**17)*1+(2**8)*229+  0, 
(2**17)*0+(2**8)* 31+ 20, (2**17)*0+(2**8)*119+121, (2**17)*0+(2**8)*122+ 91, (2**17)*0+(2**8)*128+ 83, (2**17)*0+(2**8)*144+ 70, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*230+  0, (2**17)*1+(2**8)*232+158, 
(2**17)*0+(2**8)*  6+ 50, (2**17)*0+(2**8)* 74+154, (2**17)*0+(2**8)*120+ 87, (2**17)*0+(2**8)*125+ 40, (2**17)*0+(2**8)*130+176, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*231+  0, (2**17)*1+(2**8)*236+  4, 
(2**17)*0+(2**8)* 40+102, (2**17)*0+(2**8)*123+154, (2**17)*0+(2**8)*128+ 84, (2**17)*0+(2**8)*171+157, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*215+ 97, (2**17)*0+(2**8)*221+167, (2**17)*1+(2**8)*232+  0, 
(2**17)*0+(2**8)*  6+ 61, (2**17)*0+(2**8)* 10+136, (2**17)*0+(2**8)* 43+159, (2**17)*0+(2**8)* 62+ 58, (2**17)*0+(2**8)*104+172, (2**17)*0+(2**8)*134+122, (2**17)*0+(2**8)*173+  0, (2**17)*1+(2**8)*233+  0, 
(2**17)*0+(2**8)* 70+124, (2**17)*0+(2**8)*128+ 45, (2**17)*0+(2**8)*131+162, (2**17)*0+(2**8)*137+ 33, (2**17)*0+(2**8)*169+ 74, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*200+ 61, (2**17)*1+(2**8)*234+  0, 
(2**17)*0+(2**8)*  8+ 88, (2**17)*0+(2**8)*124+119, (2**17)*0+(2**8)*140+ 17, (2**17)*0+(2**8)*152+ 55, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*226+ 92, (2**17)*0+(2**8)*235+  0, (2**17)*1+(2**8)*238+ 47, 
(2**17)*0+(2**8)*  9+  5, (2**17)*0+(2**8)* 46+133, (2**17)*0+(2**8)*122+121, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*179+ 43, (2**17)*0+(2**8)*220+ 35, (2**17)*0+(2**8)*229+ 29, (2**17)*1+(2**8)*236+  0, 
(2**17)*0+(2**8)*  3+128, (2**17)*0+(2**8)* 10+ 35, (2**17)*0+(2**8)* 43+ 91, (2**17)*0+(2**8)* 63+111, (2**17)*0+(2**8)* 83+ 83, (2**17)*0+(2**8)*169+ 43, (2**17)*0+(2**8)*177+  0, (2**17)*1+(2**8)*237+  0, 
(2**17)*0+(2**8)*  8+165, (2**17)*0+(2**8)* 89+ 20, (2**17)*0+(2**8)*124+ 25, (2**17)*0+(2**8)*125+ 81, (2**17)*0+(2**8)*172+ 32, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*187+ 78, (2**17)*1+(2**8)*238+  0, 
(2**17)*0+(2**8)*  8+122, (2**17)*0+(2**8)*110+ 11, (2**17)*0+(2**8)*121+148, (2**17)*0+(2**8)*123+ 36, (2**17)*0+(2**8)*124+  5, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*221+143, (2**17)*1+(2**8)*239+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  2+154, (2**17)*0+(2**8)* 10+ 98, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)*126+141, (2**17)*0+(2**8)*138+ 78, (2**17)*0+(2**8)*141+108, (2**17)*0+(2**8)*166+ 49, (2**17)*0+(2**8)*194+ 94, (2**17)*0+(2**8)*204+ 30, (2**17)*1+(2**8)*229+ 87, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)*  9+ 23, (2**17)*0+(2**8)* 39+159, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 62+134, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)*129+ 90, (2**17)*0+(2**8)*138+ 41, (2**17)*0+(2**8)*142+  5, (2**17)*0+(2**8)*175+ 91, (2**17)*0+(2**8)*217+105, (2**17)*1+(2**8)*248+166, 
(2**17)*0+(2**8)*  1+ 75, (2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)*  7+169, (2**17)*0+(2**8)* 30+ 35, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 51+ 88, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*114+166, (2**17)*0+(2**8)*137+136, (2**17)*0+(2**8)*175+174, (2**17)*0+(2**8)*220+164, (2**17)*1+(2**8)*225+ 79, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  5+ 70, (2**17)*0+(2**8)*  7+ 44, (2**17)*0+(2**8)*  8+  6, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 48+131, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*134+ 32, (2**17)*0+(2**8)*143+155, (2**17)*0+(2**8)*152+146, (2**17)*0+(2**8)*185+ 78, (2**17)*1+(2**8)*258+ 83, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 45+ 14, (2**17)*0+(2**8)* 46+140, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*100+ 10, (2**17)*0+(2**8)*137+161, (2**17)*0+(2**8)*145+ 79, (2**17)*0+(2**8)*146+174, (2**17)*0+(2**8)*164+ 96, (2**17)*0+(2**8)*171+ 21, (2**17)*1+(2**8)*242+ 95, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  5+139, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 73+178, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*131+168, (2**17)*0+(2**8)*140+ 16, (2**17)*0+(2**8)*144+ 81, (2**17)*0+(2**8)*165+ 39, (2**17)*0+(2**8)*167+153, (2**17)*0+(2**8)*212+135, (2**17)*1+(2**8)*229+ 16, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  8+102, (2**17)*0+(2**8)*  9+  6, (2**17)*0+(2**8)* 12+ 97, (2**17)*0+(2**8)* 16+149, (2**17)*0+(2**8)* 48+ 35, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 89+ 69, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*140+158, (2**17)*0+(2**8)*233+ 54, (2**17)*1+(2**8)*241+ 31, 
(2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)* 13+ 75, (2**17)*0+(2**8)* 19+ 80, (2**17)*0+(2**8)* 47+ 30, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*108+ 99, (2**17)*0+(2**8)*144+141, (2**17)*0+(2**8)*149+ 91, (2**17)*0+(2**8)*168+158, (2**17)*0+(2**8)*201+ 44, (2**17)*1+(2**8)*258+150, 
(2**17)*0+(2**8)*  4+ 18, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 10+112, (2**17)*0+(2**8)* 12+164, (2**17)*0+(2**8)* 21+ 49, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*116+ 73, (2**17)*0+(2**8)*143+ 40, (2**17)*0+(2**8)*190+ 20, (2**17)*0+(2**8)*224+ 86, (2**17)*1+(2**8)*231+ 86, 
(2**17)*0+(2**8)*  2+ 71, (2**17)*0+(2**8)*  4+120, (2**17)*0+(2**8)*  6+ 45, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 57+  6, (2**17)*0+(2**8)* 87+ 13, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*136+154, (2**17)*0+(2**8)*164+143, (2**17)*0+(2**8)*243+136, (2**17)*1+(2**8)*246+ 45, 
(2**17)*0+(2**8)*  1+170, (2**17)*0+(2**8)*  4+ 54, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 78+172, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*100+ 20, (2**17)*0+(2**8)*144+ 74, (2**17)*0+(2**8)*147+ 41, (2**17)*0+(2**8)*148+  6, (2**17)*0+(2**8)*198+ 90, (2**17)*1+(2**8)*234+133, 
(2**17)*0+(2**8)*  0+  9, (2**17)*0+(2**8)*  5+ 60, (2**17)*0+(2**8)*  8+ 64, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 15+133, (2**17)*0+(2**8)* 23+ 84, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 56+ 19, (2**17)*0+(2**8)* 57+138, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*122+136, (2**17)*1+(2**8)*232+ 29, 
(2**17)*0+(2**8)*  0+ 36, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 13+ 29, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*104+ 87, (2**17)*0+(2**8)*137+ 89, (2**17)*0+(2**8)*147+ 55, (2**17)*0+(2**8)*166+155, (2**17)*0+(2**8)*187+168, (2**17)*0+(2**8)*211+107, (2**17)*1+(2**8)*225+ 39, 
(2**17)*0+(2**8)*  4+103, (2**17)*0+(2**8)* 11+ 21, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 13+ 99, (2**17)*0+(2**8)* 53+ 56, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*110+140, (2**17)*0+(2**8)*145+103, (2**17)*0+(2**8)*176+125, (2**17)*0+(2**8)*203+ 20, (2**17)*1+(2**8)*242+ 52, 
(2**17)*0+(2**8)*  3+131, (2**17)*0+(2**8)* 12+177, (2**17)*0+(2**8)* 13+147, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*116+ 95, (2**17)*0+(2**8)*139+108, (2**17)*0+(2**8)*157+ 30, (2**17)*0+(2**8)*186+179, (2**17)*0+(2**8)*197+ 16, (2**17)*1+(2**8)*240+ 68, 
(2**17)*0+(2**8)* 10+ 73, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 26+ 68, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 68+ 65, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*125+ 28, (2**17)*0+(2**8)*139+ 14, (2**17)*0+(2**8)*142+134, (2**17)*0+(2**8)*153+161, (2**17)*0+(2**8)*221+171, (2**17)*1+(2**8)*237+ 40, 
(2**17)*0+(2**8)*  3+ 81, (2**17)*0+(2**8)*  6+ 98, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 85+ 94, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*114+ 79, (2**17)*0+(2**8)*141+ 52, (2**17)*0+(2**8)*144+109, (2**17)*0+(2**8)*170+ 59, (2**17)*0+(2**8)*219+ 95, (2**17)*1+(2**8)*226+ 44, 
(2**17)*0+(2**8)*  2+168, (2**17)*0+(2**8)*  3+159, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 28+ 96, (2**17)*0+(2**8)* 39+ 85, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 69+166, (2**17)*0+(2**8)* 88+ 26, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*129+113, (2**17)*0+(2**8)*138+148, (2**17)*1+(2**8)*237+126, 
(2**17)*0+(2**8)*  6+115, (2**17)*0+(2**8)*  6+114, (2**17)*0+(2**8)* 11+120, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 50+156, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*119+154, (2**17)*0+(2**8)*142+102, (2**17)*0+(2**8)*149+161, (2**17)*0+(2**8)*195+109, (2**17)*1+(2**8)*256+128, 
(2**17)*0+(2**8)*  1+126, (2**17)*0+(2**8)*  4+162, (2**17)*0+(2**8)* 13+173, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 35+167, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 77+171, (2**17)*0+(2**8)* 87+ 88, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*147+ 24, (2**17)*0+(2**8)*231+ 28, (2**17)*1+(2**8)*262+104, 
(2**17)*0+(2**8)* 10+123, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 27+ 83, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*113+ 19, (2**17)*0+(2**8)*140+155, (2**17)*0+(2**8)*143+ 10, (2**17)*0+(2**8)*173+ 68, (2**17)*0+(2**8)*181+111, (2**17)*0+(2**8)*209+ 52, (2**17)*1+(2**8)*267+161, 
(2**17)*0+(2**8)*  1+ 22, (2**17)*0+(2**8)*  2+ 70, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 56+ 90, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 82+ 53, (2**17)*0+(2**8)*110+ 49, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*139+ 85, (2**17)*0+(2**8)*146+123, (2**17)*0+(2**8)*151+ 77, (2**17)*1+(2**8)*238+166, 
(2**17)*0+(2**8)*  0+ 30, (2**17)*0+(2**8)*  2+151, (2**17)*0+(2**8)*  9+ 81, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 84+ 31, (2**17)*0+(2**8)* 98+174, (2**17)*0+(2**8)*112+  0, (2**17)*0+(2**8)*139+127, (2**17)*0+(2**8)*143+ 67, (2**17)*0+(2**8)*216+ 92, (2**17)*1+(2**8)*255+132, 
(2**17)*0+(2**8)*  0+ 58, (2**17)*0+(2**8)*  6+ 87, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 23+100, (2**17)*0+(2**8)* 36+ 12, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)*109+138, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*140+ 82, (2**17)*0+(2**8)*190+172, (2**17)*0+(2**8)*199+ 94, (2**17)*1+(2**8)*241+ 44, 
(2**17)*0+(2**8)* 11+164, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 38+107, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 78+ 97, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*135+149, (2**17)*0+(2**8)*144+ 38, (2**17)*0+(2**8)*162+162, (2**17)*0+(2**8)*215+173, (2**17)*0+(2**8)*259+146, (2**17)*1+(2**8)*268+124, 
(2**17)*0+(2**8)*  8+ 69, (2**17)*0+(2**8)*  9+ 53, (2**17)*0+(2**8)* 11+128, (2**17)*0+(2**8)* 22+155, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 79+170, (2**17)*0+(2**8)* 81+ 33, (2**17)*0+(2**8)* 92+ 85, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*118+142, (2**17)*1+(2**8)*177+152, 
(2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*120+124, (2**17)*0+(2**8)*135+ 88, (2**17)*0+(2**8)*142+136, (2**17)*0+(2**8)*149+ 34, (2**17)*0+(2**8)*149+ 73, (2**17)*0+(2**8)*160+ 81, (2**17)*0+(2**8)*193+ 79, (2**17)*0+(2**8)*202+ 43, (2**17)*1+(2**8)*263+171, 
(2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 34+146, (2**17)*0+(2**8)* 47+ 91, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*118+  3, (2**17)*0+(2**8)*141+ 89, (2**17)*0+(2**8)*143+158, (2**17)*0+(2**8)*144+ 55, (2**17)*0+(2**8)*155+ 37, (2**17)*0+(2**8)*208+ 85, (2**17)*1+(2**8)*232+ 88, 
(2**17)*0+(2**8)* 14+ 97, (2**17)*0+(2**8)* 25+ 79, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 43+ 95, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)*112+ 94, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*145+ 80, (2**17)*0+(2**8)*149+175, (2**17)*0+(2**8)*206+ 48, (2**17)*0+(2**8)*210+146, (2**17)*1+(2**8)*263+156, 
(2**17)*0+(2**8)*  5+ 63, (2**17)*0+(2**8)* 11+  1, (2**17)*0+(2**8)* 12+ 16, (2**17)*0+(2**8)* 18+ 22, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 80+ 32, (2**17)*0+(2**8)* 92+143, (2**17)*0+(2**8)*104+ 85, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*135+ 28, (2**17)*1+(2**8)*184+ 17, 
(2**17)*0+(2**8)*  3+ 17, (2**17)*0+(2**8)*  6+ 66, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*141+ 38, (2**17)*0+(2**8)*145+ 83, (2**17)*0+(2**8)*155+ 44, (2**17)*0+(2**8)*200+157, (2**17)*0+(2**8)*205+ 62, (2**17)*0+(2**8)*226+154, (2**17)*1+(2**8)*261+ 72, 
(2**17)*0+(2**8)*  0+162, (2**17)*0+(2**8)*  4+169, (2**17)*0+(2**8)*  7+ 49, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 71+140, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*134+161, (2**17)*0+(2**8)*148+ 47, (2**17)*0+(2**8)*179+ 30, (2**17)*0+(2**8)*194+ 16, (2**17)*1+(2**8)*234+116, 
(2**17)*0+(2**8)*  2+ 87, (2**17)*0+(2**8)*  3+ 42, (2**17)*0+(2**8)* 17+148, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 45+ 11, (2**17)*0+(2**8)* 70+ 70, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)*119+ 74, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*127+ 76, (2**17)*0+(2**8)*136+127, (2**17)*1+(2**8)*143+ 39, 
(2**17)*0+(2**8)* 14+124, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 42+ 69, (2**17)*0+(2**8)* 65+ 14, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)* 95+102, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*145+113, (2**17)*0+(2**8)*149+168, (2**17)*0+(2**8)*172+ 23, (2**17)*0+(2**8)*187+135, (2**17)*1+(2**8)*265+ 54, 
(2**17)*0+(2**8)*  2+149, (2**17)*0+(2**8)* 12+176, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 34+ 27, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)*105+145, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*142+ 83, (2**17)*0+(2**8)*172+ 12, (2**17)*0+(2**8)*193+ 46, (2**17)*0+(2**8)*196+126, (2**17)*1+(2**8)*244+ 64, 
(2**17)*0+(2**8)*  3+ 64, (2**17)*0+(2**8)* 11+  2, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)*122+179, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*140+ 18, (2**17)*0+(2**8)*149+143, (2**17)*0+(2**8)*161+152, (2**17)*0+(2**8)*188+ 72, (2**17)*0+(2**8)*221+ 87, (2**17)*1+(2**8)*247+154, 
(2**17)*0+(2**8)*  3+ 87, (2**17)*0+(2**8)*  5+176, (2**17)*0+(2**8)*  6+170, (2**17)*0+(2**8)* 13+ 92, (2**17)*0+(2**8)* 28+ 27, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 79+ 82, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)*117+  4, (2**17)*0+(2**8)*124+161, (2**17)*0+(2**8)*126+  0, (2**17)*1+(2**8)*201+154, 
(2**17)*0+(2**8)* 13+ 88, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 76+155, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*133+ 57, (2**17)*0+(2**8)*136+142, (2**17)*0+(2**8)*144+ 36, (2**17)*0+(2**8)*147+ 30, (2**17)*0+(2**8)*149+ 54, (2**17)*0+(2**8)*189+166, (2**17)*1+(2**8)*236+126, 
(2**17)*0+(2**8)* 10+  5, (2**17)*0+(2**8)* 21+ 69, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 64+ 32, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 88+ 96, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*142+141, (2**17)*0+(2**8)*149+152, (2**17)*0+(2**8)*168+122, (2**17)*0+(2**8)*260+125, (2**17)*1+(2**8)*265+133, 
(2**17)*0+(2**8)*  7+ 23, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*135+ 82, (2**17)*0+(2**8)*145+146, (2**17)*0+(2**8)*154+ 48, (2**17)*0+(2**8)*167+ 67, (2**17)*0+(2**8)*184+  4, (2**17)*0+(2**8)*218+ 54, (2**17)*0+(2**8)*236+103, (2**17)*1+(2**8)*246+ 15, 
(2**17)*0+(2**8)*  0+124, (2**17)*0+(2**8)* 12+ 79, (2**17)*0+(2**8)* 13+ 42, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 67+ 44, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*103+ 29, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*135+ 71, (2**17)*0+(2**8)*146+118, (2**17)*0+(2**8)*196+ 70, (2**17)*1+(2**8)*256+160, 
(2**17)*0+(2**8)*  8+ 93, (2**17)*0+(2**8)* 11+ 88, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 44+130, (2**17)*0+(2**8)* 83+123, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)* 95+ 65, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*132+ 89, (2**17)*0+(2**8)*140+105, (2**17)*0+(2**8)*148+  9, (2**17)*1+(2**8)*207+136, 
(2**17)*0+(2**8)*  1+  9, (2**17)*0+(2**8)*  3+ 97, (2**17)*0+(2**8)* 24+157, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*136+  4, (2**17)*0+(2**8)*159+ 33, (2**17)*0+(2**8)*189+141, (2**17)*0+(2**8)*198+101, (2**17)*0+(2**8)*228+ 91, (2**17)*1+(2**8)*252+ 55, 
(2**17)*0+(2**8)*  4+ 23, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 72+129, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)*115+166, (2**17)*0+(2**8)*115+ 98, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*136+ 30, (2**17)*0+(2**8)*137+ 19, (2**17)*0+(2**8)*146+ 84, (2**17)*0+(2**8)*176+ 51, (2**17)*1+(2**8)*209+157, 
(2**17)*0+(2**8)*  1+ 80, (2**17)*0+(2**8)* 43+ 87, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 60+ 84, (2**17)*0+(2**8)* 75+106, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)* 93+ 19, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*142+  7, (2**17)*0+(2**8)*147+ 57, (2**17)*0+(2**8)*150+ 35, (2**17)*1+(2**8)*266+ 68, 
(2**17)*0+(2**8)*  3+ 77, (2**17)*0+(2**8)*  6+107, (2**17)*0+(2**8)* 31+ 48, (2**17)*0+(2**8)* 59+ 93, (2**17)*0+(2**8)* 69+ 29, (2**17)*0+(2**8)* 94+ 86, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*137+154, (2**17)*0+(2**8)*145+ 98, (2**17)*0+(2**8)*180+  0, (2**17)*0+(2**8)*225+  0, (2**17)*1+(2**8)*261+141, 
(2**17)*0+(2**8)*  3+ 40, (2**17)*0+(2**8)*  7+  4, (2**17)*0+(2**8)* 40+ 90, (2**17)*0+(2**8)* 82+104, (2**17)*0+(2**8)*113+165, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*144+ 23, (2**17)*0+(2**8)*174+159, (2**17)*0+(2**8)*181+  0, (2**17)*0+(2**8)*197+134, (2**17)*0+(2**8)*226+  0, (2**17)*1+(2**8)*264+ 90, 
(2**17)*0+(2**8)*  2+135, (2**17)*0+(2**8)* 40+173, (2**17)*0+(2**8)* 85+163, (2**17)*0+(2**8)* 90+ 78, (2**17)*0+(2**8)*136+ 75, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*142+169, (2**17)*0+(2**8)*165+ 35, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*186+ 88, (2**17)*0+(2**8)*227+  0, (2**17)*1+(2**8)*249+166, 
(2**17)*0+(2**8)*  8+154, (2**17)*0+(2**8)* 17+145, (2**17)*0+(2**8)* 50+ 77, (2**17)*0+(2**8)*123+ 82, (2**17)*0+(2**8)*138+  0, (2**17)*0+(2**8)*140+ 70, (2**17)*0+(2**8)*142+ 44, (2**17)*0+(2**8)*143+  6, (2**17)*0+(2**8)*183+  0, (2**17)*0+(2**8)*183+131, (2**17)*0+(2**8)*228+  0, (2**17)*1+(2**8)*269+ 32, 
(2**17)*0+(2**8)*  2+160, (2**17)*0+(2**8)* 10+ 78, (2**17)*0+(2**8)* 11+173, (2**17)*0+(2**8)* 29+ 95, (2**17)*0+(2**8)* 36+ 20, (2**17)*0+(2**8)*107+ 94, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*180+ 14, (2**17)*0+(2**8)*181+140, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*229+  0, (2**17)*1+(2**8)*235+ 10, 
(2**17)*0+(2**8)*  5+ 15, (2**17)*0+(2**8)*  9+ 80, (2**17)*0+(2**8)* 30+ 38, (2**17)*0+(2**8)* 32+152, (2**17)*0+(2**8)* 77+134, (2**17)*0+(2**8)* 94+ 15, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*140+139, (2**17)*0+(2**8)*185+  0, (2**17)*0+(2**8)*208+178, (2**17)*0+(2**8)*230+  0, (2**17)*1+(2**8)*266+168, 
(2**17)*0+(2**8)*  5+157, (2**17)*0+(2**8)* 98+ 53, (2**17)*0+(2**8)*106+ 30, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*143+102, (2**17)*0+(2**8)*144+  6, (2**17)*0+(2**8)*147+ 97, (2**17)*0+(2**8)*151+149, (2**17)*0+(2**8)*183+ 35, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*224+ 69, (2**17)*1+(2**8)*231+  0, 
(2**17)*0+(2**8)*  9+140, (2**17)*0+(2**8)* 14+ 90, (2**17)*0+(2**8)* 33+157, (2**17)*0+(2**8)* 66+ 43, (2**17)*0+(2**8)*123+149, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*148+ 75, (2**17)*0+(2**8)*154+ 80, (2**17)*0+(2**8)*182+ 30, (2**17)*0+(2**8)*187+  0, (2**17)*0+(2**8)*232+  0, (2**17)*1+(2**8)*243+ 99, 
(2**17)*0+(2**8)*  8+ 39, (2**17)*0+(2**8)* 55+ 19, (2**17)*0+(2**8)* 89+ 85, (2**17)*0+(2**8)* 96+ 85, (2**17)*0+(2**8)*139+ 18, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*145+112, (2**17)*0+(2**8)*147+164, (2**17)*0+(2**8)*156+ 49, (2**17)*0+(2**8)*188+  0, (2**17)*0+(2**8)*233+  0, (2**17)*1+(2**8)*251+ 73, 
(2**17)*0+(2**8)*  1+153, (2**17)*0+(2**8)* 29+142, (2**17)*0+(2**8)*108+135, (2**17)*0+(2**8)*111+ 44, (2**17)*0+(2**8)*137+ 71, (2**17)*0+(2**8)*139+120, (2**17)*0+(2**8)*141+ 45, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*189+  0, (2**17)*0+(2**8)*192+  6, (2**17)*0+(2**8)*222+ 13, (2**17)*1+(2**8)*234+  0, 
(2**17)*0+(2**8)*  9+ 73, (2**17)*0+(2**8)* 12+ 40, (2**17)*0+(2**8)* 13+  5, (2**17)*0+(2**8)* 63+ 89, (2**17)*0+(2**8)* 99+132, (2**17)*0+(2**8)*136+170, (2**17)*0+(2**8)*139+ 54, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*190+  0, (2**17)*0+(2**8)*213+172, (2**17)*0+(2**8)*235+  0, (2**17)*1+(2**8)*235+ 20, 
(2**17)*0+(2**8)* 97+ 28, (2**17)*0+(2**8)*135+  9, (2**17)*0+(2**8)*140+ 60, (2**17)*0+(2**8)*143+ 64, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*150+133, (2**17)*0+(2**8)*158+ 84, (2**17)*0+(2**8)*191+  0, (2**17)*0+(2**8)*191+ 19, (2**17)*0+(2**8)*192+138, (2**17)*0+(2**8)*236+  0, (2**17)*1+(2**8)*257+136, 
(2**17)*0+(2**8)*  2+ 88, (2**17)*0+(2**8)* 12+ 54, (2**17)*0+(2**8)* 31+154, (2**17)*0+(2**8)* 52+167, (2**17)*0+(2**8)* 76+106, (2**17)*0+(2**8)* 90+ 38, (2**17)*0+(2**8)*135+ 36, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*148+ 29, (2**17)*0+(2**8)*192+  0, (2**17)*0+(2**8)*237+  0, (2**17)*1+(2**8)*239+ 87, 
(2**17)*0+(2**8)* 10+102, (2**17)*0+(2**8)* 41+124, (2**17)*0+(2**8)* 68+ 19, (2**17)*0+(2**8)*107+ 51, (2**17)*0+(2**8)*139+103, (2**17)*0+(2**8)*146+ 21, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*148+ 99, (2**17)*0+(2**8)*188+ 56, (2**17)*0+(2**8)*193+  0, (2**17)*0+(2**8)*238+  0, (2**17)*1+(2**8)*245+140, 
(2**17)*0+(2**8)*  4+107, (2**17)*0+(2**8)* 22+ 29, (2**17)*0+(2**8)* 51+178, (2**17)*0+(2**8)* 62+ 15, (2**17)*0+(2**8)*105+ 67, (2**17)*0+(2**8)*138+131, (2**17)*0+(2**8)*147+177, (2**17)*0+(2**8)*148+147, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*194+  0, (2**17)*0+(2**8)*239+  0, (2**17)*1+(2**8)*251+ 95, 
(2**17)*0+(2**8)*  4+ 13, (2**17)*0+(2**8)*  7+133, (2**17)*0+(2**8)* 18+160, (2**17)*0+(2**8)* 86+170, (2**17)*0+(2**8)*102+ 39, (2**17)*0+(2**8)*145+ 73, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*161+ 68, (2**17)*0+(2**8)*195+  0, (2**17)*0+(2**8)*203+ 65, (2**17)*0+(2**8)*240+  0, (2**17)*1+(2**8)*260+ 28, 
(2**17)*0+(2**8)*  6+ 51, (2**17)*0+(2**8)*  9+108, (2**17)*0+(2**8)* 35+ 58, (2**17)*0+(2**8)* 84+ 94, (2**17)*0+(2**8)* 91+ 43, (2**17)*0+(2**8)*138+ 81, (2**17)*0+(2**8)*141+ 98, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*220+ 94, (2**17)*0+(2**8)*241+  0, (2**17)*1+(2**8)*249+ 79, 
(2**17)*0+(2**8)*  3+147, (2**17)*0+(2**8)*102+125, (2**17)*0+(2**8)*137+168, (2**17)*0+(2**8)*138+159, (2**17)*0+(2**8)*152+  0, (2**17)*0+(2**8)*163+ 96, (2**17)*0+(2**8)*174+ 85, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*204+166, (2**17)*0+(2**8)*223+ 26, (2**17)*0+(2**8)*242+  0, (2**17)*1+(2**8)*264+113, 
(2**17)*0+(2**8)*  7+101, (2**17)*0+(2**8)* 14+160, (2**17)*0+(2**8)* 60+108, (2**17)*0+(2**8)*121+127, (2**17)*0+(2**8)*141+115, (2**17)*0+(2**8)*141+114, (2**17)*0+(2**8)*146+120, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*185+156, (2**17)*0+(2**8)*198+  0, (2**17)*0+(2**8)*243+  0, (2**17)*1+(2**8)*254+154, 
(2**17)*0+(2**8)* 12+ 23, (2**17)*0+(2**8)* 96+ 27, (2**17)*0+(2**8)*127+103, (2**17)*0+(2**8)*136+126, (2**17)*0+(2**8)*139+162, (2**17)*0+(2**8)*148+173, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*170+167, (2**17)*0+(2**8)*199+  0, (2**17)*0+(2**8)*212+171, (2**17)*0+(2**8)*222+ 88, (2**17)*1+(2**8)*244+  0, 
(2**17)*0+(2**8)*  5+154, (2**17)*0+(2**8)*  8+  9, (2**17)*0+(2**8)* 38+ 67, (2**17)*0+(2**8)* 46+110, (2**17)*0+(2**8)* 74+ 51, (2**17)*0+(2**8)*132+160, (2**17)*0+(2**8)*145+123, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*162+ 83, (2**17)*0+(2**8)*200+  0, (2**17)*0+(2**8)*245+  0, (2**17)*1+(2**8)*248+ 19, 
(2**17)*0+(2**8)*  4+ 84, (2**17)*0+(2**8)* 11+122, (2**17)*0+(2**8)* 16+ 76, (2**17)*0+(2**8)*103+165, (2**17)*0+(2**8)*136+ 22, (2**17)*0+(2**8)*137+ 70, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*191+ 90, (2**17)*0+(2**8)*201+  0, (2**17)*0+(2**8)*217+ 53, (2**17)*0+(2**8)*245+ 49, (2**17)*1+(2**8)*246+  0, 
(2**17)*0+(2**8)*  4+126, (2**17)*0+(2**8)*  8+ 66, (2**17)*0+(2**8)* 81+ 91, (2**17)*0+(2**8)*120+131, (2**17)*0+(2**8)*135+ 30, (2**17)*0+(2**8)*137+151, (2**17)*0+(2**8)*144+ 81, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*202+  0, (2**17)*0+(2**8)*219+ 31, (2**17)*0+(2**8)*233+174, (2**17)*1+(2**8)*247+  0, 
(2**17)*0+(2**8)*  5+ 81, (2**17)*0+(2**8)* 55+171, (2**17)*0+(2**8)* 64+ 93, (2**17)*0+(2**8)*106+ 43, (2**17)*0+(2**8)*135+ 58, (2**17)*0+(2**8)*141+ 87, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*158+100, (2**17)*0+(2**8)*171+ 12, (2**17)*0+(2**8)*203+  0, (2**17)*0+(2**8)*244+138, (2**17)*1+(2**8)*248+  0, 
(2**17)*0+(2**8)*  0+148, (2**17)*0+(2**8)*  9+ 37, (2**17)*0+(2**8)* 27+161, (2**17)*0+(2**8)* 80+172, (2**17)*0+(2**8)*124+145, (2**17)*0+(2**8)*133+123, (2**17)*0+(2**8)*146+164, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*173+107, (2**17)*0+(2**8)*204+  0, (2**17)*0+(2**8)*213+ 97, (2**17)*1+(2**8)*249+  0, 
(2**17)*0+(2**8)* 42+151, (2**17)*0+(2**8)*143+ 69, (2**17)*0+(2**8)*144+ 53, (2**17)*0+(2**8)*146+128, (2**17)*0+(2**8)*157+155, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*205+  0, (2**17)*0+(2**8)*214+170, (2**17)*0+(2**8)*216+ 33, (2**17)*0+(2**8)*227+ 85, (2**17)*0+(2**8)*250+  0, (2**17)*1+(2**8)*253+142, 
(2**17)*0+(2**8)*  0+ 87, (2**17)*0+(2**8)*  7+135, (2**17)*0+(2**8)* 14+ 33, (2**17)*0+(2**8)* 14+ 72, (2**17)*0+(2**8)* 25+ 80, (2**17)*0+(2**8)* 58+ 78, (2**17)*0+(2**8)* 67+ 42, (2**17)*0+(2**8)*128+170, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*206+  0, (2**17)*0+(2**8)*251+  0, (2**17)*1+(2**8)*255+124, 
(2**17)*0+(2**8)*  6+ 88, (2**17)*0+(2**8)*  8+157, (2**17)*0+(2**8)*  9+ 54, (2**17)*0+(2**8)* 20+ 36, (2**17)*0+(2**8)* 73+ 84, (2**17)*0+(2**8)* 97+ 87, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*169+146, (2**17)*0+(2**8)*182+ 91, (2**17)*0+(2**8)*207+  0, (2**17)*0+(2**8)*252+  0, (2**17)*1+(2**8)*253+  3, 
(2**17)*0+(2**8)* 10+ 79, (2**17)*0+(2**8)* 14+174, (2**17)*0+(2**8)* 71+ 47, (2**17)*0+(2**8)* 75+145, (2**17)*0+(2**8)*128+155, (2**17)*0+(2**8)*149+ 97, (2**17)*0+(2**8)*160+ 79, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*178+ 95, (2**17)*0+(2**8)*208+  0, (2**17)*0+(2**8)*247+ 94, (2**17)*1+(2**8)*253+  0, 
(2**17)*0+(2**8)*  0+ 27, (2**17)*0+(2**8)* 49+ 16, (2**17)*0+(2**8)*140+ 63, (2**17)*0+(2**8)*146+  1, (2**17)*0+(2**8)*147+ 16, (2**17)*0+(2**8)*153+ 22, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*209+  0, (2**17)*0+(2**8)*215+ 32, (2**17)*0+(2**8)*227+143, (2**17)*0+(2**8)*239+ 85, (2**17)*1+(2**8)*254+  0, 
(2**17)*0+(2**8)*  6+ 37, (2**17)*0+(2**8)* 10+ 82, (2**17)*0+(2**8)* 20+ 43, (2**17)*0+(2**8)* 65+156, (2**17)*0+(2**8)* 70+ 61, (2**17)*0+(2**8)* 91+153, (2**17)*0+(2**8)*126+ 71, (2**17)*0+(2**8)*138+ 17, (2**17)*0+(2**8)*141+ 66, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*210+  0, (2**17)*1+(2**8)*255+  0, 
(2**17)*0+(2**8)* 13+ 46, (2**17)*0+(2**8)* 44+ 29, (2**17)*0+(2**8)* 59+ 15, (2**17)*0+(2**8)* 99+115, (2**17)*0+(2**8)*135+162, (2**17)*0+(2**8)*139+169, (2**17)*0+(2**8)*142+ 49, (2**17)*0+(2**8)*166+  0, (2**17)*0+(2**8)*206+140, (2**17)*0+(2**8)*211+  0, (2**17)*0+(2**8)*256+  0, (2**17)*1+(2**8)*269+161, 
(2**17)*0+(2**8)*  1+126, (2**17)*0+(2**8)*  8+ 38, (2**17)*0+(2**8)*137+ 87, (2**17)*0+(2**8)*138+ 42, (2**17)*0+(2**8)*152+148, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*180+ 11, (2**17)*0+(2**8)*205+ 70, (2**17)*0+(2**8)*212+  0, (2**17)*0+(2**8)*254+ 74, (2**17)*0+(2**8)*257+  0, (2**17)*1+(2**8)*262+ 76, 
(2**17)*0+(2**8)* 10+112, (2**17)*0+(2**8)* 14+167, (2**17)*0+(2**8)* 37+ 22, (2**17)*0+(2**8)* 52+134, (2**17)*0+(2**8)*130+ 53, (2**17)*0+(2**8)*149+124, (2**17)*0+(2**8)*168+  0, (2**17)*0+(2**8)*177+ 69, (2**17)*0+(2**8)*200+ 14, (2**17)*0+(2**8)*213+  0, (2**17)*0+(2**8)*230+102, (2**17)*1+(2**8)*258+  0, 
(2**17)*0+(2**8)*  7+ 82, (2**17)*0+(2**8)* 37+ 11, (2**17)*0+(2**8)* 58+ 45, (2**17)*0+(2**8)* 61+125, (2**17)*0+(2**8)*109+ 63, (2**17)*0+(2**8)*137+149, (2**17)*0+(2**8)*147+176, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*169+ 27, (2**17)*0+(2**8)*214+  0, (2**17)*0+(2**8)*240+145, (2**17)*1+(2**8)*259+  0, 
(2**17)*0+(2**8)*  5+ 17, (2**17)*0+(2**8)* 14+142, (2**17)*0+(2**8)* 26+151, (2**17)*0+(2**8)* 53+ 71, (2**17)*0+(2**8)* 86+ 86, (2**17)*0+(2**8)*112+153, (2**17)*0+(2**8)*138+ 64, (2**17)*0+(2**8)*146+  2, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*215+  0, (2**17)*0+(2**8)*257+179, (2**17)*1+(2**8)*260+  0, 
(2**17)*0+(2**8)* 66+153, (2**17)*0+(2**8)*138+ 87, (2**17)*0+(2**8)*140+176, (2**17)*0+(2**8)*141+170, (2**17)*0+(2**8)*148+ 92, (2**17)*0+(2**8)*163+ 27, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*214+ 82, (2**17)*0+(2**8)*216+  0, (2**17)*0+(2**8)*252+  4, (2**17)*0+(2**8)*259+161, (2**17)*1+(2**8)*261+  0, 
(2**17)*0+(2**8)*  1+141, (2**17)*0+(2**8)*  9+ 35, (2**17)*0+(2**8)* 12+ 29, (2**17)*0+(2**8)* 14+ 53, (2**17)*0+(2**8)* 54+165, (2**17)*0+(2**8)*101+125, (2**17)*0+(2**8)*148+ 88, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*211+155, (2**17)*0+(2**8)*217+  0, (2**17)*0+(2**8)*262+  0, (2**17)*1+(2**8)*268+ 57, 
(2**17)*0+(2**8)*  7+140, (2**17)*0+(2**8)* 14+151, (2**17)*0+(2**8)* 33+121, (2**17)*0+(2**8)*125+124, (2**17)*0+(2**8)*130+132, (2**17)*0+(2**8)*145+  5, (2**17)*0+(2**8)*156+ 69, (2**17)*0+(2**8)*173+  0, (2**17)*0+(2**8)*199+ 32, (2**17)*0+(2**8)*218+  0, (2**17)*0+(2**8)*223+ 96, (2**17)*1+(2**8)*263+  0, 
(2**17)*0+(2**8)*  0+ 81, (2**17)*0+(2**8)* 10+145, (2**17)*0+(2**8)* 19+ 47, (2**17)*0+(2**8)* 32+ 66, (2**17)*0+(2**8)* 49+  3, (2**17)*0+(2**8)* 83+ 53, (2**17)*0+(2**8)*101+102, (2**17)*0+(2**8)*111+ 14, (2**17)*0+(2**8)*142+ 23, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*219+  0, (2**17)*1+(2**8)*264+  0, 
(2**17)*0+(2**8)*  0+ 70, (2**17)*0+(2**8)* 11+117, (2**17)*0+(2**8)* 61+ 69, (2**17)*0+(2**8)*121+159, (2**17)*0+(2**8)*135+124, (2**17)*0+(2**8)*147+ 79, (2**17)*0+(2**8)*148+ 42, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*202+ 44, (2**17)*0+(2**8)*220+  0, (2**17)*0+(2**8)*238+ 29, (2**17)*1+(2**8)*265+  0, 
(2**17)*0+(2**8)*  5+104, (2**17)*0+(2**8)* 13+  8, (2**17)*0+(2**8)* 72+135, (2**17)*0+(2**8)*143+ 93, (2**17)*0+(2**8)*146+ 88, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*179+130, (2**17)*0+(2**8)*218+123, (2**17)*0+(2**8)*221+  0, (2**17)*0+(2**8)*230+ 65, (2**17)*0+(2**8)*266+  0, (2**17)*1+(2**8)*267+ 89, 
(2**17)*0+(2**8)*  1+  3, (2**17)*0+(2**8)* 24+ 32, (2**17)*0+(2**8)* 54+140, (2**17)*0+(2**8)* 63+100, (2**17)*0+(2**8)* 93+ 90, (2**17)*0+(2**8)*117+ 54, (2**17)*0+(2**8)*136+  9, (2**17)*0+(2**8)*138+ 97, (2**17)*0+(2**8)*159+157, (2**17)*0+(2**8)*177+  0, (2**17)*0+(2**8)*222+  0, (2**17)*1+(2**8)*267+  0, 
(2**17)*0+(2**8)*  1+ 29, (2**17)*0+(2**8)*  2+ 18, (2**17)*0+(2**8)* 11+ 83, (2**17)*0+(2**8)* 41+ 50, (2**17)*0+(2**8)* 74+156, (2**17)*0+(2**8)*139+ 23, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*207+129, (2**17)*0+(2**8)*223+  0, (2**17)*0+(2**8)*250+166, (2**17)*0+(2**8)*250+ 98, (2**17)*1+(2**8)*268+  0, 
(2**17)*0+(2**8)*  7+  6, (2**17)*0+(2**8)* 12+ 56, (2**17)*0+(2**8)* 15+ 34, (2**17)*0+(2**8)*131+ 67, (2**17)*0+(2**8)*136+ 80, (2**17)*0+(2**8)*178+ 87, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*195+ 84, (2**17)*0+(2**8)*210+106, (2**17)*0+(2**8)*224+  0, (2**17)*0+(2**8)*228+ 19, (2**17)*1+(2**8)*269+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  6+ 52, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 49+ 36, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 81+ 17, (2**17)*0+(2**8)* 86+100, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*139+129, (2**17)*0+(2**8)*156+163, (2**17)*0+(2**8)*159+160, (2**17)*0+(2**8)*159+ 91, (2**17)*0+(2**8)*161+122, (2**17)*0+(2**8)*169+ 61, (2**17)*0+(2**8)*183+ 31, (2**17)*1+(2**8)*269+116, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 10+121, (2**17)*0+(2**8)* 14+ 48, (2**17)*0+(2**8)* 27+165, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*118+172, (2**17)*0+(2**8)*153+  4, (2**17)*0+(2**8)*161+158, (2**17)*0+(2**8)*177+145, (2**17)*0+(2**8)*185+149, (2**17)*0+(2**8)*207+ 49, (2**17)*0+(2**8)*240+ 12, (2**17)*0+(2**8)*242+180, (2**17)*1+(2**8)*265+106, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 10+109, (2**17)*0+(2**8)* 19+ 14, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 48+166, (2**17)*0+(2**8)* 67+ 29, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 78+ 78, (2**17)*0+(2**8)*106+113, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*149+ 48, (2**17)*0+(2**8)*151+ 16, (2**17)*0+(2**8)*156+ 54, (2**17)*0+(2**8)*165+171, (2**17)*0+(2**8)*262+167, (2**17)*1+(2**8)*269+ 92, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  5+ 14, (2**17)*0+(2**8)* 11+127, (2**17)*0+(2**8)* 15+ 38, (2**17)*0+(2**8)* 18+141, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 58+108, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)* 94+ 92, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*129+ 81, (2**17)*0+(2**8)*149+ 30, (2**17)*0+(2**8)*153+ 33, (2**17)*0+(2**8)*184+105, (2**17)*0+(2**8)*216+ 69, (2**17)*1+(2**8)*272+  4, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)*  6+ 13, (2**17)*0+(2**8)*  7+ 90, (2**17)*0+(2**8)* 15+ 92, (2**17)*0+(2**8)* 30+ 31, (2**17)*0+(2**8)* 31+ 88, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 49+103, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)* 84+ 45, (2**17)*0+(2**8)*112+  0, (2**17)*0+(2**8)*134+135, (2**17)*0+(2**8)*148+167, (2**17)*0+(2**8)*198+ 84, (2**17)*0+(2**8)*248+  9, (2**17)*1+(2**8)*266+  2, 
(2**17)*0+(2**8)*  0+  2, (2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 13+159, (2**17)*0+(2**8)* 22+ 61, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*129+ 86, (2**17)*0+(2**8)*149+ 57, (2**17)*0+(2**8)*153+ 63, (2**17)*0+(2**8)*160+115, (2**17)*0+(2**8)*188+112, (2**17)*0+(2**8)*195+ 10, (2**17)*0+(2**8)*241+ 31, (2**17)*0+(2**8)*249+136, (2**17)*1+(2**8)*272+  2, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  7+109, (2**17)*0+(2**8)*  8+117, (2**17)*0+(2**8)* 11+ 84, (2**17)*0+(2**8)* 27+ 35, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)* 88+171, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*132+ 76, (2**17)*0+(2**8)*135+160, (2**17)*0+(2**8)*155+ 32, (2**17)*0+(2**8)*157+ 35, (2**17)*0+(2**8)*186+ 38, (2**17)*0+(2**8)*201+ 56, (2**17)*1+(2**8)*232+ 31, 
(2**17)*0+(2**8)*  6+ 39, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)* 10+ 94, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 63+ 34, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*116+103, (2**17)*0+(2**8)*136+132, (2**17)*0+(2**8)*148+168, (2**17)*0+(2**8)*154+114, (2**17)*0+(2**8)*158+ 88, (2**17)*0+(2**8)*163+146, (2**17)*0+(2**8)*189+ 62, (2**17)*0+(2**8)*217+ 59, (2**17)*1+(2**8)*230+ 46, 
(2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)*  8+131, (2**17)*0+(2**8)* 10+124, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 52+ 18, (2**17)*0+(2**8)* 70+118, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)*112+ 48, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*144+113, (2**17)*0+(2**8)*153+ 22, (2**17)*0+(2**8)*158+ 53, (2**17)*0+(2**8)*164+124, (2**17)*0+(2**8)*221+125, (2**17)*0+(2**8)*244+ 83, (2**17)*1+(2**8)*277+ 30, 
(2**17)*0+(2**8)*  0+118, (2**17)*0+(2**8)*  1+143, (2**17)*0+(2**8)*  2+ 77, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 13+ 81, (2**17)*0+(2**8)* 26+ 99, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 60+ 55, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)*106+144, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*143+ 77, (2**17)*0+(2**8)*146+146, (2**17)*0+(2**8)*180+134, (2**17)*0+(2**8)*243+122, (2**17)*1+(2**8)*267+111, 
(2**17)*0+(2**8)*  3+ 45, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 12+ 55, (2**17)*0+(2**8)* 12+ 30, (2**17)*0+(2**8)* 13+166, (2**17)*0+(2**8)* 25+132, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 47+ 91, (2**17)*0+(2**8)* 81+123, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)* 92+143, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*120+141, (2**17)*0+(2**8)*122+ 20, (2**17)*0+(2**8)*148+ 86, (2**17)*1+(2**8)*209+ 92, 
(2**17)*0+(2**8)*  8+ 57, (2**17)*0+(2**8)*  8+119, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 12+179, (2**17)*0+(2**8)* 15+168, (2**17)*0+(2**8)* 33+162, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 90+133, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*126+125, (2**17)*0+(2**8)*136+171, (2**17)*0+(2**8)*159+  8, (2**17)*0+(2**8)*200+ 62, (2**17)*0+(2**8)*209+160, (2**17)*1+(2**8)*219+ 76, 
(2**17)*0+(2**8)*  0+178, (2**17)*0+(2**8)*  2+ 39, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 30+121, (2**17)*0+(2**8)* 46+128, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 80+123, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)* 85+ 81, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*134+ 19, (2**17)*0+(2**8)*144+  6, (2**17)*0+(2**8)*154+ 24, (2**17)*0+(2**8)*155+123, (2**17)*0+(2**8)*205+ 61, (2**17)*1+(2**8)*257+ 97, 
(2**17)*0+(2**8)*  3+  7, (2**17)*0+(2**8)*  7+ 63, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 16+ 25, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 83+ 61, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*108+101, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*148+ 72, (2**17)*0+(2**8)*153+ 79, (2**17)*0+(2**8)*173+152, (2**17)*0+(2**8)*211+134, (2**17)*0+(2**8)*214+ 26, (2**17)*0+(2**8)*220+ 45, (2**17)*1+(2**8)*275+ 49, 
(2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 15+113, (2**17)*0+(2**8)* 17+ 29, (2**17)*0+(2**8)* 22+ 98, (2**17)*0+(2**8)* 32+119, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 62+ 74, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*130+179, (2**17)*0+(2**8)*151+ 18, (2**17)*0+(2**8)*155+166, (2**17)*0+(2**8)*213+ 50, (2**17)*0+(2**8)*227+  4, (2**17)*0+(2**8)*231+157, (2**17)*1+(2**8)*271+131, 
(2**17)*0+(2**8)*  7+163, (2**17)*0+(2**8)*  7+ 56, (2**17)*0+(2**8)* 11+126, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*147+ 66, (2**17)*0+(2**8)*149+ 99, (2**17)*0+(2**8)*156+102, (2**17)*0+(2**8)*201+133, (2**17)*0+(2**8)*212+ 66, (2**17)*0+(2**8)*243+ 30, (2**17)*0+(2**8)*251+ 81, (2**17)*0+(2**8)*255+116, (2**17)*1+(2**8)*265+ 19, 
(2**17)*0+(2**8)*  6+150, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 17+ 93, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 69+ 36, (2**17)*0+(2**8)* 78+173, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*144+156, (2**17)*0+(2**8)*149+ 52, (2**17)*0+(2**8)*155+163, (2**17)*0+(2**8)*159+ 36, (2**17)*0+(2**8)*206+ 88, (2**17)*0+(2**8)*244+167, (2**17)*0+(2**8)*285+  4, (2**17)*1+(2**8)*287+ 99, 
(2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 17+ 76, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 68+ 32, (2**17)*0+(2**8)* 79+ 20, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)*124+124, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*145+ 73, (2**17)*0+(2**8)*145+ 54, (2**17)*0+(2**8)*145+ 49, (2**17)*0+(2**8)*150+161, (2**17)*0+(2**8)*152+  6, (2**17)*0+(2**8)*190+ 58, (2**17)*0+(2**8)*240+135, (2**17)*1+(2**8)*268+103, 
(2**17)*0+(2**8)*  0+139, (2**17)*0+(2**8)*  8+172, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 35+ 44, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)*104+ 99, (2**17)*0+(2**8)*126+  0, (2**17)*0+(2**8)*153+127, (2**17)*0+(2**8)*156+115, (2**17)*0+(2**8)*160+ 91, (2**17)*0+(2**8)*197+166, (2**17)*0+(2**8)*203+ 21, (2**17)*0+(2**8)*237+154, (2**17)*0+(2**8)*267+118, (2**17)*1+(2**8)*271+ 86, 
(2**17)*0+(2**8)*  2+108, (2**17)*0+(2**8)* 16+ 64, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 21+142, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 82+116, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)* 97+ 25, (2**17)*0+(2**8)*110+125, (2**17)*0+(2**8)*119+135, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*148+ 19, (2**17)*0+(2**8)*149+ 80, (2**17)*0+(2**8)*155+ 76, (2**17)*0+(2**8)*182+ 68, (2**17)*1+(2**8)*198+133, 
(2**17)*0+(2**8)*  2+168, (2**17)*0+(2**8)*  2+ 41, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 29+ 42, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*147+ 60, (2**17)*0+(2**8)*158+111, (2**17)*0+(2**8)*161+ 41, (2**17)*0+(2**8)*183+  5, (2**17)*0+(2**8)*196+ 13, (2**17)*0+(2**8)*223+ 18, (2**17)*0+(2**8)*251+106, (2**17)*0+(2**8)*261+113, (2**17)*1+(2**8)*283+ 43, 
(2**17)*0+(2**8)*  1+148, (2**17)*0+(2**8)* 14+107, (2**17)*0+(2**8)* 14+ 83, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 56+ 58, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 60+149, (2**17)*0+(2**8)* 77+  9, (2**17)*0+(2**8)* 92+167, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*157+156, (2**17)*0+(2**8)*161+173, (2**17)*0+(2**8)*170+143, (2**17)*0+(2**8)*260+ 78, (2**17)*1+(2**8)*275+ 61, 
(2**17)*0+(2**8)*  6+132, (2**17)*0+(2**8)* 16+ 84, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 43+ 83, (2**17)*0+(2**8)* 45+ 67, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 76+ 78, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*111+ 61, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*138+125, (2**17)*0+(2**8)*145+  7, (2**17)*0+(2**8)*150+160, (2**17)*0+(2**8)*160+ 52, (2**17)*0+(2**8)*160+165, (2**17)*1+(2**8)*219+ 97, 
(2**17)*0+(2**8)*  4+169, (2**17)*0+(2**8)*  7+ 72, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 61+ 48, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*101+ 44, (2**17)*0+(2**8)*113+ 28, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*137+114, (2**17)*0+(2**8)*148+ 33, (2**17)*0+(2**8)*151+160, (2**17)*0+(2**8)*151+178, (2**17)*0+(2**8)*178+ 90, (2**17)*0+(2**8)*186+ 94, (2**17)*1+(2**8)*233+ 63, 
(2**17)*0+(2**8)*  0+ 88, (2**17)*0+(2**8)*  5+153, (2**17)*0+(2**8)* 11+ 60, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 55+  4, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 74+152, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*137+ 24, (2**17)*0+(2**8)*146+  8, (2**17)*0+(2**8)*149+ 95, (2**17)*0+(2**8)*159+137, (2**17)*0+(2**8)*194+134, (2**17)*0+(2**8)*247+ 99, (2**17)*1+(2**8)*253+108, 
(2**17)*0+(2**8)*  3+140, (2**17)*0+(2**8)* 13+ 11, (2**17)*0+(2**8)* 17+166, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 28+ 27, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 95+137, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*158+ 63, (2**17)*0+(2**8)*161+109, (2**17)*0+(2**8)*208+169, (2**17)*0+(2**8)*208+103, (2**17)*0+(2**8)*246+152, (2**17)*0+(2**8)*261+ 68, (2**17)*1+(2**8)*277+ 62, 
(2**17)*0+(2**8)*  6+ 20, (2**17)*0+(2**8)* 10+114, (2**17)*0+(2**8)* 13+ 61, (2**17)*0+(2**8)* 20+142, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 40+ 92, (2**17)*0+(2**8)* 50+122, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*119+139, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*145+ 52, (2**17)*0+(2**8)*153+ 58, (2**17)*0+(2**8)*218+112, (2**17)*0+(2**8)*231+ 21, (2**17)*1+(2**8)*259+ 10, 
(2**17)*0+(2**8)*  6+156, (2**17)*0+(2**8)*  9+ 65, (2**17)*0+(2**8)* 10+123, (2**17)*0+(2**8)* 13+ 20, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 44+153, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 90+ 97, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*140+104, (2**17)*0+(2**8)*152+ 62, (2**17)*0+(2**8)*159+ 56, (2**17)*0+(2**8)*210+ 62, (2**17)*0+(2**8)*229+ 84, (2**17)*1+(2**8)*286+ 56, 
(2**17)*0+(2**8)*  3+104, (2**17)*0+(2**8)*  5+149, (2**17)*0+(2**8)* 17+106, (2**17)*0+(2**8)* 24+166, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*130+ 53, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*147+ 10, (2**17)*0+(2**8)*150+ 17, (2**17)*0+(2**8)*185+ 34, (2**17)*0+(2**8)*202+170, (2**17)*0+(2**8)*237+ 71, (2**17)*0+(2**8)*245+121, (2**17)*1+(2**8)*264+  6, 
(2**17)*0+(2**8)*  2+ 98, (2**17)*0+(2**8)* 13+  7, (2**17)*0+(2**8)* 14+ 21, (2**17)*0+(2**8)* 28+159, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 53+ 17, (2**17)*0+(2**8)* 55+105, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 89+ 13, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*142+171, (2**17)*0+(2**8)*156+132, (2**17)*0+(2**8)*160+110, (2**17)*0+(2**8)*242+ 93, (2**17)*1+(2**8)*282+  7, 
(2**17)*0+(2**8)*  1+ 69, (2**17)*0+(2**8)*  2+121, (2**17)*0+(2**8)*  8+ 31, (2**17)*0+(2**8)* 14+ 41, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 35+169, (2**17)*0+(2**8)* 47+170, (2**17)*0+(2**8)* 51+ 75, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*105+ 71, (2**17)*0+(2**8)*138+  0, (2**17)*0+(2**8)*160+171, (2**17)*0+(2**8)*238+ 96, (2**17)*0+(2**8)*256+  9, (2**17)*1+(2**8)*258+ 11, 
(2**17)*0+(2**8)*  0+ 77, (2**17)*0+(2**8)*  0+174, (2**17)*0+(2**8)* 23+170, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 34+177, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 72+ 78, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*110+171, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*152+110, (2**17)*0+(2**8)*157+ 73, (2**17)*0+(2**8)*181+ 78, (2**17)*0+(2**8)*215+ 56, (2**17)*0+(2**8)*224+ 54, (2**17)*1+(2**8)*253+151, 
(2**17)*0+(2**8)* 11+156, (2**17)*0+(2**8)* 14+132, (2**17)*0+(2**8)* 31+126, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 43+ 71, (2**17)*0+(2**8)* 48+105, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 91+ 35, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*132+120, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*141+ 37, (2**17)*0+(2**8)*145+ 43, (2**17)*0+(2**8)*152+ 98, (2**17)*0+(2**8)*168+ 95, (2**17)*1+(2**8)*226+ 83, 
(2**17)*0+(2**8)*  3+ 39, (2**17)*0+(2**8)*  4+  7, (2**17)*0+(2**8)* 12+143, (2**17)*0+(2**8)* 16+ 24, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 95+ 29, (2**17)*0+(2**8)*103+ 87, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*140+ 34, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*146+ 30, (2**17)*0+(2**8)*153+ 54, (2**17)*0+(2**8)*180+159, (2**17)*0+(2**8)*210+164, (2**17)*1+(2**8)*258+ 42, 
(2**17)*0+(2**8)* 10+110, (2**17)*0+(2**8)* 18+ 58, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 84+ 51, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*147+116, (2**17)*0+(2**8)*148+ 59, (2**17)*0+(2**8)*153+ 52, (2**17)*0+(2**8)*176+102, (2**17)*0+(2**8)*181+104, (2**17)*0+(2**8)*203+122, (2**17)*0+(2**8)*217+ 26, (2**17)*0+(2**8)*259+ 29, (2**17)*1+(2**8)*270+ 95, 
(2**17)*0+(2**8)*  3+ 37, (2**17)*0+(2**8)*  4+156, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 91+ 28, (2**17)*0+(2**8)*102+113, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*135+168, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*145+107, (2**17)*0+(2**8)*154+120, (2**17)*0+(2**8)*156+ 29, (2**17)*0+(2**8)*167+ 54, (2**17)*0+(2**8)*182+ 60, (2**17)*0+(2**8)*215+ 16, (2**17)*1+(2**8)*252+137, 
(2**17)*0+(2**8)* 12+162, (2**17)*0+(2**8)* 15+159, (2**17)*0+(2**8)* 15+ 90, (2**17)*0+(2**8)* 17+121, (2**17)*0+(2**8)* 25+ 60, (2**17)*0+(2**8)* 39+ 30, (2**17)*0+(2**8)*125+115, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*150+ 52, (2**17)*0+(2**8)*180+  0, (2**17)*0+(2**8)*193+ 36, (2**17)*0+(2**8)*216+  0, (2**17)*0+(2**8)*225+ 17, (2**17)*0+(2**8)*230+100, (2**17)*0+(2**8)*252+  0, (2**17)*1+(2**8)*283+129, 
(2**17)*0+(2**8)*  9+  3, (2**17)*0+(2**8)* 17+157, (2**17)*0+(2**8)* 33+144, (2**17)*0+(2**8)* 41+148, (2**17)*0+(2**8)* 63+ 48, (2**17)*0+(2**8)* 96+ 11, (2**17)*0+(2**8)* 98+179, (2**17)*0+(2**8)*121+105, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*154+121, (2**17)*0+(2**8)*158+ 48, (2**17)*0+(2**8)*171+165, (2**17)*0+(2**8)*181+  0, (2**17)*0+(2**8)*217+  0, (2**17)*0+(2**8)*253+  0, (2**17)*1+(2**8)*262+172, 
(2**17)*0+(2**8)*  5+ 47, (2**17)*0+(2**8)*  7+ 15, (2**17)*0+(2**8)* 12+ 53, (2**17)*0+(2**8)* 21+170, (2**17)*0+(2**8)*118+166, (2**17)*0+(2**8)*125+ 91, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*154+109, (2**17)*0+(2**8)*163+ 14, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*192+166, (2**17)*0+(2**8)*211+ 29, (2**17)*0+(2**8)*218+  0, (2**17)*0+(2**8)*222+ 78, (2**17)*0+(2**8)*250+113, (2**17)*1+(2**8)*254+  0, 
(2**17)*0+(2**8)*  5+ 29, (2**17)*0+(2**8)*  9+ 32, (2**17)*0+(2**8)* 40+104, (2**17)*0+(2**8)* 72+ 68, (2**17)*0+(2**8)*128+  3, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*149+ 14, (2**17)*0+(2**8)*155+127, (2**17)*0+(2**8)*159+ 38, (2**17)*0+(2**8)*162+141, (2**17)*0+(2**8)*183+  0, (2**17)*0+(2**8)*202+108, (2**17)*0+(2**8)*219+  0, (2**17)*0+(2**8)*238+ 92, (2**17)*0+(2**8)*255+  0, (2**17)*1+(2**8)*273+ 81, 
(2**17)*0+(2**8)*  4+166, (2**17)*0+(2**8)* 54+ 83, (2**17)*0+(2**8)*104+  8, (2**17)*0+(2**8)*122+  1, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*150+ 13, (2**17)*0+(2**8)*151+ 90, (2**17)*0+(2**8)*159+ 92, (2**17)*0+(2**8)*174+ 31, (2**17)*0+(2**8)*175+ 88, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*193+103, (2**17)*0+(2**8)*220+  0, (2**17)*0+(2**8)*228+ 45, (2**17)*0+(2**8)*256+  0, (2**17)*1+(2**8)*278+135, 
(2**17)*0+(2**8)*  5+ 56, (2**17)*0+(2**8)*  9+ 62, (2**17)*0+(2**8)* 16+114, (2**17)*0+(2**8)* 44+111, (2**17)*0+(2**8)* 51+  9, (2**17)*0+(2**8)* 97+ 30, (2**17)*0+(2**8)*105+135, (2**17)*0+(2**8)*128+  1, (2**17)*0+(2**8)*144+  2, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*157+159, (2**17)*0+(2**8)*166+ 61, (2**17)*0+(2**8)*185+  0, (2**17)*0+(2**8)*221+  0, (2**17)*0+(2**8)*257+  0, (2**17)*1+(2**8)*273+ 86, 
(2**17)*0+(2**8)* 11+ 31, (2**17)*0+(2**8)* 13+ 34, (2**17)*0+(2**8)* 42+ 37, (2**17)*0+(2**8)* 57+ 55, (2**17)*0+(2**8)* 88+ 30, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*151+109, (2**17)*0+(2**8)*152+117, (2**17)*0+(2**8)*155+ 84, (2**17)*0+(2**8)*171+ 35, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*222+  0, (2**17)*0+(2**8)*232+171, (2**17)*0+(2**8)*258+  0, (2**17)*0+(2**8)*276+ 76, (2**17)*1+(2**8)*279+160, 
(2**17)*0+(2**8)*  4+167, (2**17)*0+(2**8)* 10+113, (2**17)*0+(2**8)* 14+ 87, (2**17)*0+(2**8)* 19+145, (2**17)*0+(2**8)* 45+ 61, (2**17)*0+(2**8)* 73+ 58, (2**17)*0+(2**8)* 86+ 45, (2**17)*0+(2**8)*150+ 39, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*154+ 94, (2**17)*0+(2**8)*187+  0, (2**17)*0+(2**8)*207+ 34, (2**17)*0+(2**8)*223+  0, (2**17)*0+(2**8)*259+  0, (2**17)*0+(2**8)*260+103, (2**17)*1+(2**8)*280+132, 
(2**17)*0+(2**8)*  0+112, (2**17)*0+(2**8)*  9+ 21, (2**17)*0+(2**8)* 14+ 52, (2**17)*0+(2**8)* 20+123, (2**17)*0+(2**8)* 77+124, (2**17)*0+(2**8)*100+ 82, (2**17)*0+(2**8)*133+ 29, (2**17)*0+(2**8)*152+  0, (2**17)*0+(2**8)*152+131, (2**17)*0+(2**8)*154+124, (2**17)*0+(2**8)*188+  0, (2**17)*0+(2**8)*196+ 18, (2**17)*0+(2**8)*214+118, (2**17)*0+(2**8)*224+  0, (2**17)*0+(2**8)*256+ 48, (2**17)*1+(2**8)*260+  0, 
(2**17)*0+(2**8)*  2+145, (2**17)*0+(2**8)* 36+133, (2**17)*0+(2**8)* 99+121, (2**17)*0+(2**8)*123+110, (2**17)*0+(2**8)*144+118, (2**17)*0+(2**8)*145+143, (2**17)*0+(2**8)*146+ 77, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*157+ 81, (2**17)*0+(2**8)*170+ 99, (2**17)*0+(2**8)*189+  0, (2**17)*0+(2**8)*204+ 55, (2**17)*0+(2**8)*225+  0, (2**17)*0+(2**8)*250+144, (2**17)*0+(2**8)*261+  0, (2**17)*1+(2**8)*287+ 77, 
(2**17)*0+(2**8)*  4+ 85, (2**17)*0+(2**8)* 65+ 91, (2**17)*0+(2**8)*147+ 45, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*156+ 55, (2**17)*0+(2**8)*156+ 30, (2**17)*0+(2**8)*157+166, (2**17)*0+(2**8)*169+132, (2**17)*0+(2**8)*190+  0, (2**17)*0+(2**8)*191+ 91, (2**17)*0+(2**8)*225+123, (2**17)*0+(2**8)*226+  0, (2**17)*0+(2**8)*236+143, (2**17)*0+(2**8)*262+  0, (2**17)*0+(2**8)*264+141, (2**17)*1+(2**8)*266+ 20, 
(2**17)*0+(2**8)* 15+  7, (2**17)*0+(2**8)* 56+ 61, (2**17)*0+(2**8)* 65+159, (2**17)*0+(2**8)* 75+ 75, (2**17)*0+(2**8)*152+ 57, (2**17)*0+(2**8)*152+119, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*156+179, (2**17)*0+(2**8)*159+168, (2**17)*0+(2**8)*177+162, (2**17)*0+(2**8)*191+  0, (2**17)*0+(2**8)*227+  0, (2**17)*0+(2**8)*234+133, (2**17)*0+(2**8)*263+  0, (2**17)*0+(2**8)*270+125, (2**17)*1+(2**8)*280+171, 
(2**17)*0+(2**8)*  0+  5, (2**17)*0+(2**8)* 10+ 23, (2**17)*0+(2**8)* 11+122, (2**17)*0+(2**8)* 61+ 60, (2**17)*0+(2**8)*113+ 96, (2**17)*0+(2**8)*144+178, (2**17)*0+(2**8)*146+ 39, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*174+121, (2**17)*0+(2**8)*190+128, (2**17)*0+(2**8)*192+  0, (2**17)*0+(2**8)*224+123, (2**17)*0+(2**8)*228+  0, (2**17)*0+(2**8)*229+ 81, (2**17)*0+(2**8)*264+  0, (2**17)*1+(2**8)*278+ 19, 
(2**17)*0+(2**8)*  4+ 71, (2**17)*0+(2**8)*  9+ 78, (2**17)*0+(2**8)* 29+151, (2**17)*0+(2**8)* 67+133, (2**17)*0+(2**8)* 70+ 25, (2**17)*0+(2**8)* 76+ 44, (2**17)*0+(2**8)*131+ 48, (2**17)*0+(2**8)*147+  7, (2**17)*0+(2**8)*151+ 63, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*160+ 25, (2**17)*0+(2**8)*193+  0, (2**17)*0+(2**8)*227+ 61, (2**17)*0+(2**8)*229+  0, (2**17)*0+(2**8)*252+101, (2**17)*1+(2**8)*265+  0, 
(2**17)*0+(2**8)*  7+ 17, (2**17)*0+(2**8)* 11+165, (2**17)*0+(2**8)* 69+ 49, (2**17)*0+(2**8)* 83+  3, (2**17)*0+(2**8)* 87+156, (2**17)*0+(2**8)*127+130, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*159+113, (2**17)*0+(2**8)*161+ 29, (2**17)*0+(2**8)*166+ 98, (2**17)*0+(2**8)*176+119, (2**17)*0+(2**8)*194+  0, (2**17)*0+(2**8)*206+ 74, (2**17)*0+(2**8)*230+  0, (2**17)*0+(2**8)*266+  0, (2**17)*1+(2**8)*274+179, 
(2**17)*0+(2**8)*  3+ 65, (2**17)*0+(2**8)*  5+ 98, (2**17)*0+(2**8)* 12+101, (2**17)*0+(2**8)* 57+132, (2**17)*0+(2**8)* 68+ 65, (2**17)*0+(2**8)* 99+ 29, (2**17)*0+(2**8)*107+ 80, (2**17)*0+(2**8)*111+115, (2**17)*0+(2**8)*121+ 18, (2**17)*0+(2**8)*151+163, (2**17)*0+(2**8)*151+ 56, (2**17)*0+(2**8)*155+126, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*195+  0, (2**17)*0+(2**8)*231+  0, (2**17)*1+(2**8)*267+  0, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)*  5+ 51, (2**17)*0+(2**8)* 11+162, (2**17)*0+(2**8)* 15+ 35, (2**17)*0+(2**8)* 62+ 87, (2**17)*0+(2**8)*100+166, (2**17)*0+(2**8)*141+  3, (2**17)*0+(2**8)*143+ 98, (2**17)*0+(2**8)*150+150, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*161+ 93, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*213+ 36, (2**17)*0+(2**8)*222+173, (2**17)*0+(2**8)*232+  0, (2**17)*1+(2**8)*268+  0, 
(2**17)*0+(2**8)*  1+ 72, (2**17)*0+(2**8)*  1+ 53, (2**17)*0+(2**8)*  1+ 48, (2**17)*0+(2**8)*  6+160, (2**17)*0+(2**8)*  8+  5, (2**17)*0+(2**8)* 46+ 57, (2**17)*0+(2**8)* 96+134, (2**17)*0+(2**8)*124+102, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*161+ 76, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*212+ 32, (2**17)*0+(2**8)*223+ 20, (2**17)*0+(2**8)*233+  0, (2**17)*0+(2**8)*268+124, (2**17)*1+(2**8)*269+  0, 
(2**17)*0+(2**8)*  9+126, (2**17)*0+(2**8)* 12+114, (2**17)*0+(2**8)* 16+ 90, (2**17)*0+(2**8)* 53+165, (2**17)*0+(2**8)* 59+ 20, (2**17)*0+(2**8)* 93+153, (2**17)*0+(2**8)*123+117, (2**17)*0+(2**8)*127+ 85, (2**17)*0+(2**8)*144+139, (2**17)*0+(2**8)*152+172, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*179+ 44, (2**17)*0+(2**8)*198+  0, (2**17)*0+(2**8)*234+  0, (2**17)*0+(2**8)*248+ 99, (2**17)*1+(2**8)*270+  0, 
(2**17)*0+(2**8)*  4+ 18, (2**17)*0+(2**8)*  5+ 79, (2**17)*0+(2**8)* 11+ 75, (2**17)*0+(2**8)* 38+ 67, (2**17)*0+(2**8)* 54+132, (2**17)*0+(2**8)*146+108, (2**17)*0+(2**8)*160+ 64, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*165+142, (2**17)*0+(2**8)*199+  0, (2**17)*0+(2**8)*226+116, (2**17)*0+(2**8)*235+  0, (2**17)*0+(2**8)*241+ 25, (2**17)*0+(2**8)*254+125, (2**17)*0+(2**8)*263+135, (2**17)*1+(2**8)*271+  0, 
(2**17)*0+(2**8)*  3+ 59, (2**17)*0+(2**8)* 14+110, (2**17)*0+(2**8)* 17+ 40, (2**17)*0+(2**8)* 39+  4, (2**17)*0+(2**8)* 52+ 12, (2**17)*0+(2**8)* 79+ 17, (2**17)*0+(2**8)*107+105, (2**17)*0+(2**8)*117+112, (2**17)*0+(2**8)*139+ 42, (2**17)*0+(2**8)*146+168, (2**17)*0+(2**8)*146+ 41, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*173+ 42, (2**17)*0+(2**8)*200+  0, (2**17)*0+(2**8)*236+  0, (2**17)*1+(2**8)*272+  0, 
(2**17)*0+(2**8)* 13+155, (2**17)*0+(2**8)* 17+172, (2**17)*0+(2**8)* 26+142, (2**17)*0+(2**8)*116+ 77, (2**17)*0+(2**8)*131+ 60, (2**17)*0+(2**8)*145+148, (2**17)*0+(2**8)*158+107, (2**17)*0+(2**8)*158+ 83, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*200+ 58, (2**17)*0+(2**8)*201+  0, (2**17)*0+(2**8)*204+149, (2**17)*0+(2**8)*221+  9, (2**17)*0+(2**8)*236+167, (2**17)*0+(2**8)*237+  0, (2**17)*1+(2**8)*273+  0, 
(2**17)*0+(2**8)*  1+  6, (2**17)*0+(2**8)*  6+159, (2**17)*0+(2**8)* 16+ 51, (2**17)*0+(2**8)* 16+164, (2**17)*0+(2**8)* 75+ 96, (2**17)*0+(2**8)*150+132, (2**17)*0+(2**8)*160+ 84, (2**17)*0+(2**8)*166+  0, (2**17)*0+(2**8)*187+ 83, (2**17)*0+(2**8)*189+ 67, (2**17)*0+(2**8)*202+  0, (2**17)*0+(2**8)*220+ 78, (2**17)*0+(2**8)*238+  0, (2**17)*0+(2**8)*255+ 61, (2**17)*0+(2**8)*274+  0, (2**17)*1+(2**8)*282+125, 
(2**17)*0+(2**8)*  4+ 32, (2**17)*0+(2**8)*  7+159, (2**17)*0+(2**8)*  7+177, (2**17)*0+(2**8)* 34+ 89, (2**17)*0+(2**8)* 42+ 93, (2**17)*0+(2**8)* 89+ 62, (2**17)*0+(2**8)*148+169, (2**17)*0+(2**8)*151+ 72, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*203+  0, (2**17)*0+(2**8)*205+ 48, (2**17)*0+(2**8)*239+  0, (2**17)*0+(2**8)*245+ 44, (2**17)*0+(2**8)*257+ 28, (2**17)*0+(2**8)*275+  0, (2**17)*1+(2**8)*281+114, 
(2**17)*0+(2**8)*  2+  7, (2**17)*0+(2**8)*  5+ 94, (2**17)*0+(2**8)* 15+136, (2**17)*0+(2**8)* 50+133, (2**17)*0+(2**8)*103+ 98, (2**17)*0+(2**8)*109+107, (2**17)*0+(2**8)*144+ 88, (2**17)*0+(2**8)*149+153, (2**17)*0+(2**8)*155+ 60, (2**17)*0+(2**8)*168+  0, (2**17)*0+(2**8)*199+  4, (2**17)*0+(2**8)*204+  0, (2**17)*0+(2**8)*218+152, (2**17)*0+(2**8)*240+  0, (2**17)*0+(2**8)*276+  0, (2**17)*1+(2**8)*281+ 24, 
(2**17)*0+(2**8)* 14+ 62, (2**17)*0+(2**8)* 17+108, (2**17)*0+(2**8)* 64+168, (2**17)*0+(2**8)* 64+102, (2**17)*0+(2**8)*102+151, (2**17)*0+(2**8)*117+ 67, (2**17)*0+(2**8)*133+ 61, (2**17)*0+(2**8)*147+140, (2**17)*0+(2**8)*157+ 11, (2**17)*0+(2**8)*161+166, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*172+ 27, (2**17)*0+(2**8)*205+  0, (2**17)*0+(2**8)*239+137, (2**17)*0+(2**8)*241+  0, (2**17)*1+(2**8)*277+  0, 
(2**17)*0+(2**8)*  1+ 51, (2**17)*0+(2**8)*  9+ 57, (2**17)*0+(2**8)* 74+111, (2**17)*0+(2**8)* 87+ 20, (2**17)*0+(2**8)*115+  9, (2**17)*0+(2**8)*150+ 20, (2**17)*0+(2**8)*154+114, (2**17)*0+(2**8)*157+ 61, (2**17)*0+(2**8)*164+142, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*184+ 92, (2**17)*0+(2**8)*194+122, (2**17)*0+(2**8)*206+  0, (2**17)*0+(2**8)*242+  0, (2**17)*0+(2**8)*263+139, (2**17)*1+(2**8)*278+  0, 
(2**17)*0+(2**8)*  8+ 61, (2**17)*0+(2**8)* 15+ 55, (2**17)*0+(2**8)* 66+ 61, (2**17)*0+(2**8)* 85+ 83, (2**17)*0+(2**8)*142+ 55, (2**17)*0+(2**8)*150+156, (2**17)*0+(2**8)*153+ 65, (2**17)*0+(2**8)*154+123, (2**17)*0+(2**8)*157+ 20, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*188+153, (2**17)*0+(2**8)*207+  0, (2**17)*0+(2**8)*234+ 97, (2**17)*0+(2**8)*243+  0, (2**17)*0+(2**8)*279+  0, (2**17)*1+(2**8)*284+104, 
(2**17)*0+(2**8)*  3+  9, (2**17)*0+(2**8)*  6+ 16, (2**17)*0+(2**8)* 41+ 33, (2**17)*0+(2**8)* 58+169, (2**17)*0+(2**8)* 93+ 70, (2**17)*0+(2**8)*101+120, (2**17)*0+(2**8)*120+  5, (2**17)*0+(2**8)*147+104, (2**17)*0+(2**8)*149+149, (2**17)*0+(2**8)*161+106, (2**17)*0+(2**8)*168+166, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*208+  0, (2**17)*0+(2**8)*244+  0, (2**17)*0+(2**8)*274+ 53, (2**17)*1+(2**8)*280+  0, 
(2**17)*0+(2**8)* 12+131, (2**17)*0+(2**8)* 16+109, (2**17)*0+(2**8)* 98+ 92, (2**17)*0+(2**8)*138+  6, (2**17)*0+(2**8)*146+ 98, (2**17)*0+(2**8)*157+  7, (2**17)*0+(2**8)*158+ 21, (2**17)*0+(2**8)*172+159, (2**17)*0+(2**8)*173+  0, (2**17)*0+(2**8)*197+ 17, (2**17)*0+(2**8)*199+105, (2**17)*0+(2**8)*209+  0, (2**17)*0+(2**8)*233+ 13, (2**17)*0+(2**8)*245+  0, (2**17)*0+(2**8)*281+  0, (2**17)*1+(2**8)*286+171, 
(2**17)*0+(2**8)* 16+170, (2**17)*0+(2**8)* 94+ 95, (2**17)*0+(2**8)*112+  8, (2**17)*0+(2**8)*114+ 10, (2**17)*0+(2**8)*145+ 69, (2**17)*0+(2**8)*146+121, (2**17)*0+(2**8)*152+ 31, (2**17)*0+(2**8)*158+ 41, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*179+169, (2**17)*0+(2**8)*191+170, (2**17)*0+(2**8)*195+ 75, (2**17)*0+(2**8)*210+  0, (2**17)*0+(2**8)*246+  0, (2**17)*0+(2**8)*249+ 71, (2**17)*1+(2**8)*282+  0, 
(2**17)*0+(2**8)*  8+109, (2**17)*0+(2**8)* 13+ 72, (2**17)*0+(2**8)* 37+ 77, (2**17)*0+(2**8)* 71+ 55, (2**17)*0+(2**8)* 80+ 53, (2**17)*0+(2**8)*109+150, (2**17)*0+(2**8)*144+ 77, (2**17)*0+(2**8)*144+174, (2**17)*0+(2**8)*167+170, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*178+177, (2**17)*0+(2**8)*211+  0, (2**17)*0+(2**8)*216+ 78, (2**17)*0+(2**8)*247+  0, (2**17)*0+(2**8)*254+171, (2**17)*1+(2**8)*283+  0, 
(2**17)*0+(2**8)*  1+ 42, (2**17)*0+(2**8)*  8+ 97, (2**17)*0+(2**8)* 24+ 94, (2**17)*0+(2**8)* 82+ 82, (2**17)*0+(2**8)*155+156, (2**17)*0+(2**8)*158+132, (2**17)*0+(2**8)*175+126, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*187+ 71, (2**17)*0+(2**8)*192+105, (2**17)*0+(2**8)*212+  0, (2**17)*0+(2**8)*235+ 35, (2**17)*0+(2**8)*248+  0, (2**17)*0+(2**8)*276+120, (2**17)*0+(2**8)*284+  0, (2**17)*1+(2**8)*285+ 37, 
(2**17)*0+(2**8)*  2+ 29, (2**17)*0+(2**8)*  9+ 53, (2**17)*0+(2**8)* 36+158, (2**17)*0+(2**8)* 66+163, (2**17)*0+(2**8)*114+ 41, (2**17)*0+(2**8)*147+ 39, (2**17)*0+(2**8)*148+  7, (2**17)*0+(2**8)*156+143, (2**17)*0+(2**8)*160+ 24, (2**17)*0+(2**8)*177+  0, (2**17)*0+(2**8)*213+  0, (2**17)*0+(2**8)*239+ 29, (2**17)*0+(2**8)*247+ 87, (2**17)*0+(2**8)*249+  0, (2**17)*0+(2**8)*284+ 34, (2**17)*1+(2**8)*285+  0, 
(2**17)*0+(2**8)*  3+115, (2**17)*0+(2**8)*  4+ 58, (2**17)*0+(2**8)*  9+ 51, (2**17)*0+(2**8)* 32+101, (2**17)*0+(2**8)* 37+103, (2**17)*0+(2**8)* 59+121, (2**17)*0+(2**8)* 73+ 25, (2**17)*0+(2**8)*115+ 28, (2**17)*0+(2**8)*126+ 94, (2**17)*0+(2**8)*154+110, (2**17)*0+(2**8)*162+ 58, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*214+  0, (2**17)*0+(2**8)*228+ 51, (2**17)*0+(2**8)*250+  0, (2**17)*1+(2**8)*286+  0, 
(2**17)*0+(2**8)*  1+106, (2**17)*0+(2**8)* 10+119, (2**17)*0+(2**8)* 12+ 28, (2**17)*0+(2**8)* 23+ 53, (2**17)*0+(2**8)* 38+ 59, (2**17)*0+(2**8)* 71+ 15, (2**17)*0+(2**8)*108+136, (2**17)*0+(2**8)*147+ 37, (2**17)*0+(2**8)*148+156, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*215+  0, (2**17)*0+(2**8)*235+ 28, (2**17)*0+(2**8)*246+113, (2**17)*0+(2**8)*251+  0, (2**17)*0+(2**8)*279+168, (2**17)*1+(2**8)*287+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  3+156, (2**17)*0+(2**8)*  6+166, (2**17)*0+(2**8)*  8+ 43, (2**17)*0+(2**8)*  9+ 64, (2**17)*0+(2**8)* 13+ 71, (2**17)*0+(2**8)* 14+ 60, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 40+ 44, (2**17)*0+(2**8)* 54+140, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 72+140, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)* 97+ 54, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*164+ 10, (2**17)*0+(2**8)*228+ 11, (2**17)*0+(2**8)*268+ 81, (2**17)*0+(2**8)*286+ 56, (2**17)*1+(2**8)*290+ 76, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)* 15+127, (2**17)*0+(2**8)* 19+142, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 31+ 44, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)*101+102, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*151+101, (2**17)*0+(2**8)*152+ 52, (2**17)*0+(2**8)*152+ 95, (2**17)*0+(2**8)*157+132, (2**17)*0+(2**8)*163+112, (2**17)*0+(2**8)*196+137, (2**17)*0+(2**8)*217+ 86, (2**17)*0+(2**8)*219+106, (2**17)*0+(2**8)*250+ 96, (2**17)*0+(2**8)*281+ 22, (2**17)*1+(2**8)*298+ 36, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 12+159, (2**17)*0+(2**8)* 28+ 59, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 42+ 93, (2**17)*0+(2**8)* 56+ 84, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 70+111, (2**17)*0+(2**8)* 91+ 60, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)*116+  6, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*130+102, (2**17)*0+(2**8)*150+ 49, (2**17)*0+(2**8)*155+ 68, (2**17)*0+(2**8)*159+110, (2**17)*0+(2**8)*162+123, (2**17)*0+(2**8)*177+ 85, (2**17)*0+(2**8)*215+ 78, (2**17)*1+(2**8)*282+177, 
(2**17)*0+(2**8)*  0+112, (2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  4+164, (2**17)*0+(2**8)*  8+ 48, (2**17)*0+(2**8)* 12+177, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 34+125, (2**17)*0+(2**8)* 58+120, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 79+  6, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*137+176, (2**17)*0+(2**8)*148+ 78, (2**17)*0+(2**8)*155+ 62, (2**17)*0+(2**8)*161+177, (2**17)*0+(2**8)*167+122, (2**17)*0+(2**8)*214+109, (2**17)*0+(2**8)*240+ 53, (2**17)*1+(2**8)*261+ 13, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)*  5+119, (2**17)*0+(2**8)*  8+ 17, (2**17)*0+(2**8)* 15+105, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 39+ 66, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 87+101, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*109+151, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*137+ 71, (2**17)*0+(2**8)*146+107, (2**17)*0+(2**8)*154+131, (2**17)*0+(2**8)*159+ 35, (2**17)*0+(2**8)*159+ 52, (2**17)*0+(2**8)*161+  7, (2**17)*0+(2**8)*205+  7, (2**17)*0+(2**8)*227+ 48, (2**17)*1+(2**8)*263+ 44, 
(2**17)*0+(2**8)*  2+ 83, (2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)*  7+ 79, (2**17)*0+(2**8)* 12+ 12, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 48+ 55, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 89+ 48, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*132+149, (2**17)*0+(2**8)*152+170, (2**17)*0+(2**8)*154+ 81, (2**17)*0+(2**8)*158+ 37, (2**17)*0+(2**8)*163+ 63, (2**17)*0+(2**8)*205+138, (2**17)*0+(2**8)*213+177, (2**17)*0+(2**8)*241+ 68, (2**17)*0+(2**8)*265+ 35, (2**17)*1+(2**8)*297+ 63, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  9+ 63, (2**17)*0+(2**8)* 17+113, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 45+ 75, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*111+122, (2**17)*0+(2**8)*126+  0, (2**17)*0+(2**8)*129+161, (2**17)*0+(2**8)*143+ 35, (2**17)*0+(2**8)*150+ 54, (2**17)*0+(2**8)*153+167, (2**17)*0+(2**8)*156+139, (2**17)*0+(2**8)*157+ 70, (2**17)*0+(2**8)*161+ 61, (2**17)*0+(2**8)*187+155, (2**17)*0+(2**8)*223+153, (2**17)*0+(2**8)*236+ 76, (2**17)*1+(2**8)*257+134, 
(2**17)*0+(2**8)*  2+121, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  7+ 26, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 62+  1, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 83+ 96, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*116+ 78, (2**17)*0+(2**8)*123+ 61, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*151+107, (2**17)*0+(2**8)*153+ 72, (2**17)*0+(2**8)*157+ 29, (2**17)*0+(2**8)*172+159, (2**17)*0+(2**8)*177+ 18, (2**17)*0+(2**8)*197+103, (2**17)*0+(2**8)*202+ 19, (2**17)*0+(2**8)*242+ 29, (2**17)*1+(2**8)*270+131, 
(2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 12+126, (2**17)*0+(2**8)* 22+171, (2**17)*0+(2**8)* 28+132, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*100+131, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*130+118, (2**17)*0+(2**8)*151+150, (2**17)*0+(2**8)*153+168, (2**17)*0+(2**8)*153+ 86, (2**17)*0+(2**8)*163+147, (2**17)*0+(2**8)*189+  6, (2**17)*0+(2**8)*206+106, (2**17)*0+(2**8)*212+121, (2**17)*0+(2**8)*221+171, (2**17)*0+(2**8)*244+132, (2**17)*1+(2**8)*291+114, 
(2**17)*0+(2**8)*  2+150, (2**17)*0+(2**8)*  8+ 28, (2**17)*0+(2**8)*  8+ 74, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 58+ 33, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 77+141, (2**17)*0+(2**8)* 82+151, (2**17)*0+(2**8)* 98+158, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*105+ 50, (2**17)*0+(2**8)*121+ 28, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*133+ 60, (2**17)*0+(2**8)*154+ 40, (2**17)*0+(2**8)*156+ 87, (2**17)*0+(2**8)*156+ 12, (2**17)*0+(2**8)*163+124, (2**17)*1+(2**8)*203+ 94, 
(2**17)*0+(2**8)*  3+ 56, (2**17)*0+(2**8)*  4+ 51, (2**17)*0+(2**8)*  9+ 24, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 18+ 99, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 76+ 28, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*128+ 55, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*150+ 43, (2**17)*0+(2**8)*164+109, (2**17)*0+(2**8)*174+ 93, (2**17)*0+(2**8)*184+157, (2**17)*0+(2**8)*199+ 26, (2**17)*0+(2**8)*233+ 68, (2**17)*0+(2**8)*253+ 10, (2**17)*0+(2**8)*267+166, (2**17)*1+(2**8)*283+119, 
(2**17)*0+(2**8)*  1+ 50, (2**17)*0+(2**8)*  5+131, (2**17)*0+(2**8)*  6+172, (2**17)*0+(2**8)*  6+ 33, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 12+ 42, (2**17)*0+(2**8)* 13+119, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 45+ 58, (2**17)*0+(2**8)* 63+147, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 89+ 34, (2**17)*0+(2**8)* 90+178, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*115+ 10, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*145+ 36, (2**17)*0+(2**8)*161+143, (2**17)*0+(2**8)*209+ 30, (2**17)*1+(2**8)*294+115, 
(2**17)*0+(2**8)*  2+ 68, (2**17)*0+(2**8)*  7+179, (2**17)*0+(2**8)*  9+ 25, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 37+ 28, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 86+148, (2**17)*0+(2**8)* 98+111, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*102+152, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*135+134, (2**17)*0+(2**8)*150+ 73, (2**17)*0+(2**8)*160+158, (2**17)*0+(2**8)*161+ 65, (2**17)*0+(2**8)*179+ 63, (2**17)*0+(2**8)*196+ 70, (2**17)*0+(2**8)*231+112, (2**17)*1+(2**8)*296+ 68, 
(2**17)*0+(2**8)*  0+143, (2**17)*0+(2**8)*  1+155, (2**17)*0+(2**8)*  4+139, (2**17)*0+(2**8)*  9+143, (2**17)*0+(2**8)* 12+ 27, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)* 87+ 14, (2**17)*0+(2**8)* 88+ 98, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*157+115, (2**17)*0+(2**8)*163+138, (2**17)*0+(2**8)*192+ 95, (2**17)*0+(2**8)*193+159, (2**17)*0+(2**8)*252+ 81, (2**17)*0+(2**8)*269+ 23, (2**17)*0+(2**8)*292+ 57, (2**17)*1+(2**8)*294+ 65, 
(2**17)*0+(2**8)*  3+  7, (2**17)*0+(2**8)* 12+  1, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 32+ 46, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 59+ 86, (2**17)*0+(2**8)* 61+ 70, (2**17)*0+(2**8)* 71+160, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*155+ 35, (2**17)*0+(2**8)*156+ 22, (2**17)*0+(2**8)*157+163, (2**17)*0+(2**8)*159+ 91, (2**17)*0+(2**8)*161+137, (2**17)*0+(2**8)*263+131, (2**17)*0+(2**8)*267+145, (2**17)*0+(2**8)*275+ 71, (2**17)*1+(2**8)*277+ 66, 
(2**17)*0+(2**8)*  5+ 57, (2**17)*0+(2**8)* 10+166, (2**17)*0+(2**8)* 11+132, (2**17)*0+(2**8)* 14+ 33, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 25+  9, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 51+111, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*106+  3, (2**17)*0+(2**8)*108+153, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*136+ 48, (2**17)*0+(2**8)*150+107, (2**17)*0+(2**8)*155+110, (2**17)*0+(2**8)*181+161, (2**17)*0+(2**8)*222+134, (2**17)*0+(2**8)*230+ 69, (2**17)*1+(2**8)*276+171, 
(2**17)*0+(2**8)*  0+ 69, (2**17)*0+(2**8)*  2+145, (2**17)*0+(2**8)*  5+ 31, (2**17)*0+(2**8)*  8+108, (2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 36+174, (2**17)*0+(2**8)* 43+ 15, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 61+ 56, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*108+ 25, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*138+108, (2**17)*0+(2**8)*151+ 30, (2**17)*0+(2**8)*164+ 91, (2**17)*0+(2**8)*179+ 54, (2**17)*0+(2**8)*232+154, (2**17)*0+(2**8)*264+ 11, (2**17)*1+(2**8)*279+106, 
(2**17)*0+(2**8)*  1+ 49, (2**17)*0+(2**8)*  1+170, (2**17)*0+(2**8)*  2+ 46, (2**17)*0+(2**8)*  6+ 65, (2**17)*0+(2**8)*  9+ 84, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 38+167, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)* 95+ 10, (2**17)*0+(2**8)* 99+124, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*154+ 39, (2**17)*0+(2**8)*176+ 64, (2**17)*0+(2**8)*190+ 85, (2**17)*0+(2**8)*219+ 92, (2**17)*0+(2**8)*224+118, (2**17)*0+(2**8)*289+147, (2**17)*1+(2**8)*299+134, 
(2**17)*0+(2**8)* 11+166, (2**17)*0+(2**8)* 16+108, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 38+ 67, (2**17)*0+(2**8)* 41+ 14, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 67+131, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*119+117, (2**17)*0+(2**8)*123+165, (2**17)*0+(2**8)*138+  0, (2**17)*0+(2**8)*153+ 19, (2**17)*0+(2**8)*155+  6, (2**17)*0+(2**8)*157+ 65, (2**17)*0+(2**8)*160+ 31, (2**17)*0+(2**8)*164+ 13, (2**17)*0+(2**8)*230+117, (2**17)*0+(2**8)*255+ 38, (2**17)*1+(2**8)*284+153, 
(2**17)*0+(2**8)*  1+ 41, (2**17)*0+(2**8)*  1+ 72, (2**17)*0+(2**8)* 10+106, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 57+ 85, (2**17)*0+(2**8)* 60+ 59, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)* 94+ 32, (2**17)*0+(2**8)*106+ 40, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*122+ 39, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*140+ 33, (2**17)*0+(2**8)*150+ 83, (2**17)*0+(2**8)*152+165, (2**17)*0+(2**8)*157+167, (2**17)*0+(2**8)*173+156, (2**17)*0+(2**8)*201+ 68, (2**17)*1+(2**8)*216+ 24, 
(2**17)*0+(2**8)*  5+172, (2**17)*0+(2**8)*  5+ 46, (2**17)*0+(2**8)*  8+ 90, (2**17)*0+(2**8)* 14+  3, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 26+143, (2**17)*0+(2**8)* 30+ 40, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 65+ 88, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*124+115, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*155+ 98, (2**17)*0+(2**8)*171+ 20, (2**17)*0+(2**8)*185+ 31, (2**17)*0+(2**8)*223+ 94, (2**17)*0+(2**8)*249+ 53, (2**17)*0+(2**8)*254+155, (2**17)*1+(2**8)*272+168, 
(2**17)*0+(2**8)*  9+ 55, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 23+ 36, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 64+ 20, (2**17)*0+(2**8)* 70+ 82, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*121+ 63, (2**17)*0+(2**8)*126+130, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*154+122, (2**17)*0+(2**8)*156+ 52, (2**17)*0+(2**8)*156+ 27, (2**17)*0+(2**8)*158+  2, (2**17)*0+(2**8)*164+113, (2**17)*0+(2**8)*183+ 89, (2**17)*0+(2**8)*183+ 34, (2**17)*0+(2**8)*253+160, (2**17)*1+(2**8)*262+105, 
(2**17)*0+(2**8)* 13+ 41, (2**17)*0+(2**8)* 14+148, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)*109+134, (2**17)*0+(2**8)*112+  0, (2**17)*0+(2**8)*141+153, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*150+ 52, (2**17)*0+(2**8)*153+151, (2**17)*0+(2**8)*159+165, (2**17)*0+(2**8)*160+173, (2**17)*0+(2**8)*163+ 35, (2**17)*0+(2**8)*182+ 41, (2**17)*0+(2**8)*197+170, (2**17)*0+(2**8)*231+ 27, (2**17)*0+(2**8)*235+ 93, (2**17)*0+(2**8)*251+179, (2**17)*1+(2**8)*284+152, 
(2**17)*0+(2**8)*  8+100, (2**17)*0+(2**8)* 13+ 83, (2**17)*0+(2**8)* 13+153, (2**17)*0+(2**8)* 14+ 18, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 54+141, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 84+ 62, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*114+ 38, (2**17)*0+(2**8)*135+103, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*143+150, (2**17)*0+(2**8)*160+122, (2**17)*0+(2**8)*169+ 30, (2**17)*0+(2**8)*171+163, (2**17)*0+(2**8)*191+ 58, (2**17)*0+(2**8)*229+ 91, (2**17)*1+(2**8)*262+ 64, 
(2**17)*0+(2**8)*  1+ 91, (2**17)*0+(2**8)*  3+ 65, (2**17)*0+(2**8)*  4+ 13, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 60+ 24, (2**17)*0+(2**8)* 68+171, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)* 96+142, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*152+148, (2**17)*0+(2**8)*157+ 77, (2**17)*0+(2**8)*170+103, (2**17)*0+(2**8)*170+131, (2**17)*0+(2**8)*186+163, (2**17)*0+(2**8)*207+103, (2**17)*0+(2**8)*246+ 23, (2**17)*0+(2**8)*274+ 32, (2**17)*1+(2**8)*292+ 29, 
(2**17)*0+(2**8)*  3+169, (2**17)*0+(2**8)* 10+ 76, (2**17)*0+(2**8)* 13+168, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 30+117, (2**17)*0+(2**8)* 53+ 51, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*118+ 34, (2**17)*0+(2**8)*139+127, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*153+ 80, (2**17)*0+(2**8)*161+ 40, (2**17)*0+(2**8)*162+130, (2**17)*0+(2**8)*162+152, (2**17)*0+(2**8)*218+ 74, (2**17)*0+(2**8)*225+ 57, (2**17)*0+(2**8)*260+ 35, (2**17)*1+(2**8)*295+ 65, 
(2**17)*0+(2**8)* 10+ 29, (2**17)*0+(2**8)* 10+ 93, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 50+ 79, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 76+ 64, (2**17)*0+(2**8)* 78+103, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)* 95+  3, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*150+  7, (2**17)*0+(2**8)*156+ 58, (2**17)*0+(2**8)*160+109, (2**17)*0+(2**8)*160+ 41, (2**17)*0+(2**8)*175+ 26, (2**17)*0+(2**8)*202+ 17, (2**17)*0+(2**8)*247+178, (2**17)*0+(2**8)*288+176, (2**17)*1+(2**8)*297+159, 
(2**17)*0+(2**8)*  4+119, (2**17)*0+(2**8)*  8+176, (2**17)*0+(2**8)* 11+154, (2**17)*0+(2**8)* 12+114, (2**17)*0+(2**8)* 14+ 75, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 44+ 68, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 75+150, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*104+104, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*131+130, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*149+122, (2**17)*0+(2**8)*157+ 54, (2**17)*0+(2**8)*162+107, (2**17)*0+(2**8)*200+ 45, (2**17)*0+(2**8)*234+154, (2**17)*1+(2**8)*257+ 26, 
(2**17)*0+(2**8)*  1+121, (2**17)*0+(2**8)*  4+ 25, (2**17)*0+(2**8)*  8+ 49, (2**17)*0+(2**8)* 10+142, (2**17)*0+(2**8)* 11+ 99, (2**17)*0+(2**8)* 18+ 28, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 48+ 94, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)* 92+  5, (2**17)*0+(2**8)*110+149, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*127+127, (2**17)*0+(2**8)*128+ 91, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*164+162, (2**17)*0+(2**8)*185+ 39, (2**17)*0+(2**8)*224+148, (2**17)*1+(2**8)*235+117, 
(2**17)*0+(2**8)*  0+148, (2**17)*0+(2**8)*  2+ 36, (2**17)*0+(2**8)*  4+  5, (2**17)*0+(2**8)* 11+121, (2**17)*0+(2**8)* 16+153, (2**17)*0+(2**8)* 24+ 32, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 49+ 57, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 66+162, (2**17)*0+(2**8)* 88+134, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*120+ 29, (2**17)*0+(2**8)*125+ 94, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*156+ 99, (2**17)*0+(2**8)*194+ 26, (2**17)*0+(2**8)*243+ 37, (2**17)*1+(2**8)*243+155, 
(2**17)*0+(2**8)* 14+  9, (2**17)*0+(2**8)* 78+ 10, (2**17)*0+(2**8)*118+ 80, (2**17)*0+(2**8)*136+ 55, (2**17)*0+(2**8)*140+ 75, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*153+156, (2**17)*0+(2**8)*156+166, (2**17)*0+(2**8)*158+ 43, (2**17)*0+(2**8)*159+ 64, (2**17)*0+(2**8)*163+ 71, (2**17)*0+(2**8)*164+ 60, (2**17)*0+(2**8)*180+  0, (2**17)*0+(2**8)*190+ 44, (2**17)*0+(2**8)*204+140, (2**17)*0+(2**8)*210+  0, (2**17)*0+(2**8)*222+140, (2**17)*0+(2**8)*240+  0, (2**17)*0+(2**8)*247+ 54, (2**17)*1+(2**8)*270+  0, 
(2**17)*0+(2**8)*  1+100, (2**17)*0+(2**8)*  2+ 51, (2**17)*0+(2**8)*  2+ 94, (2**17)*0+(2**8)*  7+131, (2**17)*0+(2**8)* 13+111, (2**17)*0+(2**8)* 46+136, (2**17)*0+(2**8)* 67+ 85, (2**17)*0+(2**8)* 69+105, (2**17)*0+(2**8)*100+ 95, (2**17)*0+(2**8)*131+ 21, (2**17)*0+(2**8)*148+ 35, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*165+127, (2**17)*0+(2**8)*169+142, (2**17)*0+(2**8)*181+  0, (2**17)*0+(2**8)*181+ 44, (2**17)*0+(2**8)*211+  0, (2**17)*0+(2**8)*241+  0, (2**17)*0+(2**8)*251+102, (2**17)*1+(2**8)*271+  0, 
(2**17)*0+(2**8)*  0+ 48, (2**17)*0+(2**8)*  5+ 67, (2**17)*0+(2**8)*  9+109, (2**17)*0+(2**8)* 12+122, (2**17)*0+(2**8)* 27+ 84, (2**17)*0+(2**8)* 65+ 77, (2**17)*0+(2**8)*132+176, (2**17)*0+(2**8)*152+  0, (2**17)*0+(2**8)*162+159, (2**17)*0+(2**8)*178+ 59, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*192+ 93, (2**17)*0+(2**8)*206+ 84, (2**17)*0+(2**8)*212+  0, (2**17)*0+(2**8)*220+111, (2**17)*0+(2**8)*241+ 60, (2**17)*0+(2**8)*242+  0, (2**17)*0+(2**8)*266+  6, (2**17)*0+(2**8)*272+  0, (2**17)*1+(2**8)*280+102, 
(2**17)*0+(2**8)*  5+ 61, (2**17)*0+(2**8)* 11+176, (2**17)*0+(2**8)* 17+121, (2**17)*0+(2**8)* 64+108, (2**17)*0+(2**8)* 90+ 52, (2**17)*0+(2**8)*111+ 12, (2**17)*0+(2**8)*150+112, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*154+164, (2**17)*0+(2**8)*158+ 48, (2**17)*0+(2**8)*162+177, (2**17)*0+(2**8)*183+  0, (2**17)*0+(2**8)*184+125, (2**17)*0+(2**8)*208+120, (2**17)*0+(2**8)*213+  0, (2**17)*0+(2**8)*229+  6, (2**17)*0+(2**8)*243+  0, (2**17)*0+(2**8)*273+  0, (2**17)*0+(2**8)*287+176, (2**17)*1+(2**8)*298+ 78, 
(2**17)*0+(2**8)*  4+130, (2**17)*0+(2**8)*  9+ 34, (2**17)*0+(2**8)*  9+ 51, (2**17)*0+(2**8)* 11+  6, (2**17)*0+(2**8)* 55+  6, (2**17)*0+(2**8)* 77+ 47, (2**17)*0+(2**8)*113+ 43, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*155+119, (2**17)*0+(2**8)*158+ 17, (2**17)*0+(2**8)*165+105, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*189+ 66, (2**17)*0+(2**8)*214+  0, (2**17)*0+(2**8)*237+101, (2**17)*0+(2**8)*244+  0, (2**17)*0+(2**8)*259+151, (2**17)*0+(2**8)*274+  0, (2**17)*0+(2**8)*287+ 71, (2**17)*1+(2**8)*296+107, 
(2**17)*0+(2**8)*  2+169, (2**17)*0+(2**8)*  4+ 80, (2**17)*0+(2**8)*  8+ 36, (2**17)*0+(2**8)* 13+ 62, (2**17)*0+(2**8)* 55+137, (2**17)*0+(2**8)* 63+176, (2**17)*0+(2**8)* 91+ 67, (2**17)*0+(2**8)*115+ 34, (2**17)*0+(2**8)*147+ 62, (2**17)*0+(2**8)*152+ 83, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*157+ 79, (2**17)*0+(2**8)*162+ 12, (2**17)*0+(2**8)*185+  0, (2**17)*0+(2**8)*198+ 55, (2**17)*0+(2**8)*215+  0, (2**17)*0+(2**8)*239+ 48, (2**17)*0+(2**8)*245+  0, (2**17)*0+(2**8)*275+  0, (2**17)*1+(2**8)*282+149, 
(2**17)*0+(2**8)*  0+ 53, (2**17)*0+(2**8)*  3+166, (2**17)*0+(2**8)*  6+138, (2**17)*0+(2**8)*  7+ 69, (2**17)*0+(2**8)* 11+ 60, (2**17)*0+(2**8)* 37+154, (2**17)*0+(2**8)* 73+152, (2**17)*0+(2**8)* 86+ 75, (2**17)*0+(2**8)*107+133, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*159+ 63, (2**17)*0+(2**8)*167+113, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*195+ 75, (2**17)*0+(2**8)*216+  0, (2**17)*0+(2**8)*246+  0, (2**17)*0+(2**8)*261+122, (2**17)*0+(2**8)*276+  0, (2**17)*0+(2**8)*279+161, (2**17)*1+(2**8)*293+ 35, 
(2**17)*0+(2**8)*  1+106, (2**17)*0+(2**8)*  3+ 71, (2**17)*0+(2**8)*  7+ 28, (2**17)*0+(2**8)* 22+158, (2**17)*0+(2**8)* 27+ 17, (2**17)*0+(2**8)* 47+102, (2**17)*0+(2**8)* 52+ 18, (2**17)*0+(2**8)* 92+ 28, (2**17)*0+(2**8)*120+130, (2**17)*0+(2**8)*152+121, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*157+ 26, (2**17)*0+(2**8)*187+  0, (2**17)*0+(2**8)*212+  1, (2**17)*0+(2**8)*217+  0, (2**17)*0+(2**8)*233+ 96, (2**17)*0+(2**8)*247+  0, (2**17)*0+(2**8)*266+ 78, (2**17)*0+(2**8)*273+ 61, (2**17)*1+(2**8)*277+  0, 
(2**17)*0+(2**8)*  1+149, (2**17)*0+(2**8)*  3+167, (2**17)*0+(2**8)*  3+ 85, (2**17)*0+(2**8)* 13+146, (2**17)*0+(2**8)* 39+  5, (2**17)*0+(2**8)* 56+105, (2**17)*0+(2**8)* 62+120, (2**17)*0+(2**8)* 71+170, (2**17)*0+(2**8)* 94+131, (2**17)*0+(2**8)*141+113, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*162+126, (2**17)*0+(2**8)*172+171, (2**17)*0+(2**8)*178+132, (2**17)*0+(2**8)*188+  0, (2**17)*0+(2**8)*218+  0, (2**17)*0+(2**8)*248+  0, (2**17)*0+(2**8)*250+131, (2**17)*0+(2**8)*278+  0, (2**17)*1+(2**8)*280+118, 
(2**17)*0+(2**8)*  4+ 39, (2**17)*0+(2**8)*  6+ 86, (2**17)*0+(2**8)*  6+ 11, (2**17)*0+(2**8)* 13+123, (2**17)*0+(2**8)* 53+ 93, (2**17)*0+(2**8)*152+150, (2**17)*0+(2**8)*158+ 28, (2**17)*0+(2**8)*158+ 74, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*189+  0, (2**17)*0+(2**8)*208+ 33, (2**17)*0+(2**8)*219+  0, (2**17)*0+(2**8)*227+141, (2**17)*0+(2**8)*232+151, (2**17)*0+(2**8)*248+158, (2**17)*0+(2**8)*249+  0, (2**17)*0+(2**8)*255+ 50, (2**17)*0+(2**8)*271+ 28, (2**17)*0+(2**8)*279+  0, (2**17)*1+(2**8)*283+ 60, 
(2**17)*0+(2**8)*  0+ 42, (2**17)*0+(2**8)* 14+108, (2**17)*0+(2**8)* 24+ 92, (2**17)*0+(2**8)* 34+156, (2**17)*0+(2**8)* 49+ 25, (2**17)*0+(2**8)* 83+ 67, (2**17)*0+(2**8)*103+  9, (2**17)*0+(2**8)*117+165, (2**17)*0+(2**8)*133+118, (2**17)*0+(2**8)*153+ 56, (2**17)*0+(2**8)*154+ 51, (2**17)*0+(2**8)*159+ 24, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*168+ 99, (2**17)*0+(2**8)*190+  0, (2**17)*0+(2**8)*220+  0, (2**17)*0+(2**8)*226+ 28, (2**17)*0+(2**8)*250+  0, (2**17)*0+(2**8)*278+ 55, (2**17)*1+(2**8)*280+  0, 
(2**17)*0+(2**8)* 11+142, (2**17)*0+(2**8)* 59+ 29, (2**17)*0+(2**8)*144+114, (2**17)*0+(2**8)*151+ 50, (2**17)*0+(2**8)*155+131, (2**17)*0+(2**8)*156+172, (2**17)*0+(2**8)*156+ 33, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*162+ 42, (2**17)*0+(2**8)*163+119, (2**17)*0+(2**8)*191+  0, (2**17)*0+(2**8)*195+ 58, (2**17)*0+(2**8)*213+147, (2**17)*0+(2**8)*221+  0, (2**17)*0+(2**8)*239+ 34, (2**17)*0+(2**8)*240+178, (2**17)*0+(2**8)*251+  0, (2**17)*0+(2**8)*265+ 10, (2**17)*0+(2**8)*281+  0, (2**17)*1+(2**8)*295+ 36, 
(2**17)*0+(2**8)*  0+ 72, (2**17)*0+(2**8)* 10+157, (2**17)*0+(2**8)* 11+ 64, (2**17)*0+(2**8)* 29+ 62, (2**17)*0+(2**8)* 46+ 69, (2**17)*0+(2**8)* 81+111, (2**17)*0+(2**8)*146+ 67, (2**17)*0+(2**8)*152+ 68, (2**17)*0+(2**8)*157+179, (2**17)*0+(2**8)*159+ 25, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*187+ 28, (2**17)*0+(2**8)*192+  0, (2**17)*0+(2**8)*222+  0, (2**17)*0+(2**8)*236+148, (2**17)*0+(2**8)*248+111, (2**17)*0+(2**8)*252+  0, (2**17)*0+(2**8)*252+152, (2**17)*0+(2**8)*282+  0, (2**17)*1+(2**8)*285+134, 
(2**17)*0+(2**8)*  7+114, (2**17)*0+(2**8)* 13+137, (2**17)*0+(2**8)* 42+ 94, (2**17)*0+(2**8)* 43+158, (2**17)*0+(2**8)*102+ 80, (2**17)*0+(2**8)*119+ 22, (2**17)*0+(2**8)*142+ 56, (2**17)*0+(2**8)*144+ 64, (2**17)*0+(2**8)*150+143, (2**17)*0+(2**8)*151+155, (2**17)*0+(2**8)*154+139, (2**17)*0+(2**8)*159+143, (2**17)*0+(2**8)*162+ 27, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*193+  0, (2**17)*0+(2**8)*223+  0, (2**17)*0+(2**8)*237+ 14, (2**17)*0+(2**8)*238+ 98, (2**17)*0+(2**8)*253+  0, (2**17)*1+(2**8)*283+  0, 
(2**17)*0+(2**8)*  5+ 34, (2**17)*0+(2**8)*  6+ 21, (2**17)*0+(2**8)*  7+162, (2**17)*0+(2**8)*  9+ 90, (2**17)*0+(2**8)* 11+136, (2**17)*0+(2**8)*113+130, (2**17)*0+(2**8)*117+144, (2**17)*0+(2**8)*125+ 70, (2**17)*0+(2**8)*127+ 65, (2**17)*0+(2**8)*153+  7, (2**17)*0+(2**8)*162+  1, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*182+ 46, (2**17)*0+(2**8)*194+  0, (2**17)*0+(2**8)*209+ 86, (2**17)*0+(2**8)*211+ 70, (2**17)*0+(2**8)*221+160, (2**17)*0+(2**8)*224+  0, (2**17)*0+(2**8)*254+  0, (2**17)*1+(2**8)*284+  0, 
(2**17)*0+(2**8)*  0+106, (2**17)*0+(2**8)*  5+109, (2**17)*0+(2**8)* 31+160, (2**17)*0+(2**8)* 72+133, (2**17)*0+(2**8)* 80+ 68, (2**17)*0+(2**8)*126+170, (2**17)*0+(2**8)*155+ 57, (2**17)*0+(2**8)*160+166, (2**17)*0+(2**8)*161+132, (2**17)*0+(2**8)*164+ 33, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*175+  9, (2**17)*0+(2**8)*195+  0, (2**17)*0+(2**8)*201+111, (2**17)*0+(2**8)*225+  0, (2**17)*0+(2**8)*255+  0, (2**17)*0+(2**8)*256+  3, (2**17)*0+(2**8)*258+153, (2**17)*0+(2**8)*285+  0, (2**17)*1+(2**8)*286+ 48, 
(2**17)*0+(2**8)*  1+ 29, (2**17)*0+(2**8)* 14+ 90, (2**17)*0+(2**8)* 29+ 53, (2**17)*0+(2**8)* 82+153, (2**17)*0+(2**8)*114+ 10, (2**17)*0+(2**8)*129+105, (2**17)*0+(2**8)*150+ 69, (2**17)*0+(2**8)*152+145, (2**17)*0+(2**8)*155+ 31, (2**17)*0+(2**8)*158+108, (2**17)*0+(2**8)*166+  0, (2**17)*0+(2**8)*186+174, (2**17)*0+(2**8)*193+ 15, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*211+ 56, (2**17)*0+(2**8)*226+  0, (2**17)*0+(2**8)*256+  0, (2**17)*0+(2**8)*258+ 25, (2**17)*0+(2**8)*286+  0, (2**17)*1+(2**8)*288+108, 
(2**17)*0+(2**8)*  4+ 38, (2**17)*0+(2**8)* 26+ 63, (2**17)*0+(2**8)* 40+ 84, (2**17)*0+(2**8)* 69+ 91, (2**17)*0+(2**8)* 74+117, (2**17)*0+(2**8)*139+146, (2**17)*0+(2**8)*149+133, (2**17)*0+(2**8)*151+ 49, (2**17)*0+(2**8)*151+170, (2**17)*0+(2**8)*152+ 46, (2**17)*0+(2**8)*156+ 65, (2**17)*0+(2**8)*159+ 84, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*188+167, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*227+  0, (2**17)*0+(2**8)*245+ 10, (2**17)*0+(2**8)*249+124, (2**17)*0+(2**8)*257+  0, (2**17)*1+(2**8)*287+  0, 
(2**17)*0+(2**8)*  3+ 18, (2**17)*0+(2**8)*  5+  5, (2**17)*0+(2**8)*  7+ 64, (2**17)*0+(2**8)* 10+ 30, (2**17)*0+(2**8)* 14+ 12, (2**17)*0+(2**8)* 80+116, (2**17)*0+(2**8)*105+ 37, (2**17)*0+(2**8)*134+152, (2**17)*0+(2**8)*161+166, (2**17)*0+(2**8)*166+108, (2**17)*0+(2**8)*168+  0, (2**17)*0+(2**8)*188+ 67, (2**17)*0+(2**8)*191+ 14, (2**17)*0+(2**8)*198+  0, (2**17)*0+(2**8)*217+131, (2**17)*0+(2**8)*228+  0, (2**17)*0+(2**8)*258+  0, (2**17)*0+(2**8)*269+117, (2**17)*0+(2**8)*273+165, (2**17)*1+(2**8)*288+  0, 
(2**17)*0+(2**8)*  0+ 82, (2**17)*0+(2**8)*  2+164, (2**17)*0+(2**8)*  7+166, (2**17)*0+(2**8)* 23+155, (2**17)*0+(2**8)* 51+ 67, (2**17)*0+(2**8)* 66+ 23, (2**17)*0+(2**8)*151+ 41, (2**17)*0+(2**8)*151+ 72, (2**17)*0+(2**8)*160+106, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*199+  0, (2**17)*0+(2**8)*207+ 85, (2**17)*0+(2**8)*210+ 59, (2**17)*0+(2**8)*229+  0, (2**17)*0+(2**8)*244+ 32, (2**17)*0+(2**8)*256+ 40, (2**17)*0+(2**8)*259+  0, (2**17)*0+(2**8)*272+ 39, (2**17)*0+(2**8)*289+  0, (2**17)*1+(2**8)*290+ 33, 
(2**17)*0+(2**8)*  5+ 97, (2**17)*0+(2**8)* 21+ 19, (2**17)*0+(2**8)* 35+ 30, (2**17)*0+(2**8)* 73+ 93, (2**17)*0+(2**8)* 99+ 52, (2**17)*0+(2**8)*104+154, (2**17)*0+(2**8)*122+167, (2**17)*0+(2**8)*155+172, (2**17)*0+(2**8)*155+ 46, (2**17)*0+(2**8)*158+ 90, (2**17)*0+(2**8)*164+  3, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*176+143, (2**17)*0+(2**8)*180+ 40, (2**17)*0+(2**8)*200+  0, (2**17)*0+(2**8)*215+ 88, (2**17)*0+(2**8)*230+  0, (2**17)*0+(2**8)*260+  0, (2**17)*0+(2**8)*274+115, (2**17)*1+(2**8)*290+  0, 
(2**17)*0+(2**8)*  4+121, (2**17)*0+(2**8)*  6+ 51, (2**17)*0+(2**8)*  6+ 26, (2**17)*0+(2**8)*  8+  1, (2**17)*0+(2**8)* 14+112, (2**17)*0+(2**8)* 33+ 88, (2**17)*0+(2**8)* 33+ 33, (2**17)*0+(2**8)*103+159, (2**17)*0+(2**8)*112+104, (2**17)*0+(2**8)*159+ 55, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*173+ 36, (2**17)*0+(2**8)*201+  0, (2**17)*0+(2**8)*214+ 20, (2**17)*0+(2**8)*220+ 82, (2**17)*0+(2**8)*231+  0, (2**17)*0+(2**8)*261+  0, (2**17)*0+(2**8)*271+ 63, (2**17)*0+(2**8)*276+130, (2**17)*1+(2**8)*291+  0, 
(2**17)*0+(2**8)*  0+ 51, (2**17)*0+(2**8)*  3+150, (2**17)*0+(2**8)*  9+164, (2**17)*0+(2**8)* 10+172, (2**17)*0+(2**8)* 13+ 34, (2**17)*0+(2**8)* 32+ 40, (2**17)*0+(2**8)* 47+169, (2**17)*0+(2**8)* 81+ 26, (2**17)*0+(2**8)* 85+ 92, (2**17)*0+(2**8)*101+178, (2**17)*0+(2**8)*134+151, (2**17)*0+(2**8)*163+ 41, (2**17)*0+(2**8)*164+148, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*202+  0, (2**17)*0+(2**8)*232+  0, (2**17)*0+(2**8)*259+134, (2**17)*0+(2**8)*262+  0, (2**17)*0+(2**8)*291+153, (2**17)*1+(2**8)*292+  0, 
(2**17)*0+(2**8)* 10+121, (2**17)*0+(2**8)* 19+ 29, (2**17)*0+(2**8)* 21+162, (2**17)*0+(2**8)* 41+ 57, (2**17)*0+(2**8)* 79+ 90, (2**17)*0+(2**8)*112+ 63, (2**17)*0+(2**8)*158+100, (2**17)*0+(2**8)*163+ 83, (2**17)*0+(2**8)*163+153, (2**17)*0+(2**8)*164+ 18, (2**17)*0+(2**8)*173+  0, (2**17)*0+(2**8)*203+  0, (2**17)*0+(2**8)*204+141, (2**17)*0+(2**8)*233+  0, (2**17)*0+(2**8)*234+ 62, (2**17)*0+(2**8)*263+  0, (2**17)*0+(2**8)*264+ 38, (2**17)*0+(2**8)*285+103, (2**17)*0+(2**8)*293+  0, (2**17)*1+(2**8)*293+150, 
(2**17)*0+(2**8)*  2+147, (2**17)*0+(2**8)*  7+ 76, (2**17)*0+(2**8)* 20+102, (2**17)*0+(2**8)* 20+130, (2**17)*0+(2**8)* 36+162, (2**17)*0+(2**8)* 57+102, (2**17)*0+(2**8)* 96+ 22, (2**17)*0+(2**8)*124+ 31, (2**17)*0+(2**8)*142+ 28, (2**17)*0+(2**8)*151+ 91, (2**17)*0+(2**8)*153+ 65, (2**17)*0+(2**8)*154+ 13, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*204+  0, (2**17)*0+(2**8)*210+ 24, (2**17)*0+(2**8)*218+171, (2**17)*0+(2**8)*234+  0, (2**17)*0+(2**8)*246+142, (2**17)*0+(2**8)*264+  0, (2**17)*1+(2**8)*294+  0, 
(2**17)*0+(2**8)*  3+ 79, (2**17)*0+(2**8)* 11+ 39, (2**17)*0+(2**8)* 12+129, (2**17)*0+(2**8)* 12+151, (2**17)*0+(2**8)* 68+ 73, (2**17)*0+(2**8)* 75+ 56, (2**17)*0+(2**8)*110+ 34, (2**17)*0+(2**8)*145+ 64, (2**17)*0+(2**8)*153+169, (2**17)*0+(2**8)*160+ 76, (2**17)*0+(2**8)*163+168, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*180+117, (2**17)*0+(2**8)*203+ 51, (2**17)*0+(2**8)*205+  0, (2**17)*0+(2**8)*235+  0, (2**17)*0+(2**8)*265+  0, (2**17)*0+(2**8)*268+ 34, (2**17)*0+(2**8)*289+127, (2**17)*1+(2**8)*295+  0, 
(2**17)*0+(2**8)*  0+  6, (2**17)*0+(2**8)*  6+ 57, (2**17)*0+(2**8)* 10+108, (2**17)*0+(2**8)* 10+ 40, (2**17)*0+(2**8)* 25+ 25, (2**17)*0+(2**8)* 52+ 16, (2**17)*0+(2**8)* 97+177, (2**17)*0+(2**8)*138+175, (2**17)*0+(2**8)*147+158, (2**17)*0+(2**8)*160+ 29, (2**17)*0+(2**8)*160+ 93, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*200+ 79, (2**17)*0+(2**8)*206+  0, (2**17)*0+(2**8)*226+ 64, (2**17)*0+(2**8)*228+103, (2**17)*0+(2**8)*236+  0, (2**17)*0+(2**8)*245+  3, (2**17)*0+(2**8)*266+  0, (2**17)*1+(2**8)*296+  0, 
(2**17)*0+(2**8)*  7+ 53, (2**17)*0+(2**8)* 12+106, (2**17)*0+(2**8)* 50+ 44, (2**17)*0+(2**8)* 84+153, (2**17)*0+(2**8)*107+ 25, (2**17)*0+(2**8)*154+119, (2**17)*0+(2**8)*158+176, (2**17)*0+(2**8)*161+154, (2**17)*0+(2**8)*162+114, (2**17)*0+(2**8)*164+ 75, (2**17)*0+(2**8)*177+  0, (2**17)*0+(2**8)*194+ 68, (2**17)*0+(2**8)*207+  0, (2**17)*0+(2**8)*225+150, (2**17)*0+(2**8)*237+  0, (2**17)*0+(2**8)*254+104, (2**17)*0+(2**8)*267+  0, (2**17)*0+(2**8)*281+130, (2**17)*0+(2**8)*297+  0, (2**17)*1+(2**8)*299+122, 
(2**17)*0+(2**8)* 14+161, (2**17)*0+(2**8)* 35+ 38, (2**17)*0+(2**8)* 74+147, (2**17)*0+(2**8)* 85+116, (2**17)*0+(2**8)*151+121, (2**17)*0+(2**8)*154+ 25, (2**17)*0+(2**8)*158+ 49, (2**17)*0+(2**8)*160+142, (2**17)*0+(2**8)*161+ 99, (2**17)*0+(2**8)*168+ 28, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*198+ 94, (2**17)*0+(2**8)*208+  0, (2**17)*0+(2**8)*238+  0, (2**17)*0+(2**8)*242+  5, (2**17)*0+(2**8)*260+149, (2**17)*0+(2**8)*268+  0, (2**17)*0+(2**8)*277+127, (2**17)*0+(2**8)*278+ 91, (2**17)*1+(2**8)*298+  0, 
(2**17)*0+(2**8)*  6+ 98, (2**17)*0+(2**8)* 44+ 25, (2**17)*0+(2**8)* 93+ 36, (2**17)*0+(2**8)* 93+154, (2**17)*0+(2**8)*150+148, (2**17)*0+(2**8)*152+ 36, (2**17)*0+(2**8)*154+  5, (2**17)*0+(2**8)*161+121, (2**17)*0+(2**8)*166+153, (2**17)*0+(2**8)*174+ 32, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*199+ 57, (2**17)*0+(2**8)*209+  0, (2**17)*0+(2**8)*216+162, (2**17)*0+(2**8)*238+134, (2**17)*0+(2**8)*239+  0, (2**17)*0+(2**8)*269+  0, (2**17)*0+(2**8)*270+ 29, (2**17)*0+(2**8)*275+ 94, (2**17)*1+(2**8)*299+  0, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  1+145, (2**17)*0+(2**8)* 15+ 98, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 25+156, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 57+119, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 77+ 15, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)* 83+ 11, (2**17)*0+(2**8)* 91+168, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*109+103, (2**17)*0+(2**8)*109+107, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*121+174, (2**17)*0+(2**8)*136+108, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*152+ 40, (2**17)*0+(2**8)*153+ 17, (2**17)*0+(2**8)*177+116, (2**17)*0+(2**8)*194+ 61, (2**17)*0+(2**8)*210+ 19, (2**17)*1+(2**8)*239+ 32, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)*  3+174, (2**17)*0+(2**8)*  8+ 94, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 30+164, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 43+ 40, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)* 86+ 37, (2**17)*0+(2**8)* 92+113, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*108+ 56, (2**17)*0+(2**8)*115+165, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*136+153, (2**17)*0+(2**8)*137+ 99, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*154+ 45, (2**17)*0+(2**8)*156+ 42, (2**17)*0+(2**8)*177+ 60, (2**17)*0+(2**8)*195+ 25, (2**17)*0+(2**8)*219+154, (2**17)*0+(2**8)*223+ 27, (2**17)*1+(2**8)*226+146, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 17+ 37, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 38+ 95, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 76+121, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)* 98+ 44, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*105+ 59, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*148+130, (2**17)*0+(2**8)*149+118, (2**17)*0+(2**8)*160+ 81, (2**17)*0+(2**8)*167+159, (2**17)*0+(2**8)*189+131, (2**17)*0+(2**8)*203+141, (2**17)*0+(2**8)*215+118, (2**17)*0+(2**8)*232+175, (2**17)*0+(2**8)*251+ 91, (2**17)*0+(2**8)*261+ 52, (2**17)*0+(2**8)*282+177, (2**17)*1+(2**8)*288+ 62, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  5+ 92, (2**17)*0+(2**8)* 13+148, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 36+104, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 53+ 56, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)* 90+100, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*114+ 35, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*131+156, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*145+101, (2**17)*0+(2**8)*173+ 34, (2**17)*0+(2**8)*186+ 59, (2**17)*0+(2**8)*205+145, (2**17)*0+(2**8)*223+ 87, (2**17)*0+(2**8)*239+123, (2**17)*0+(2**8)*242+ 15, (2**17)*0+(2**8)*275+130, (2**17)*0+(2**8)*294+ 87, (2**17)*1+(2**8)*316+ 62, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 16+ 41, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 44+ 13, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 74+124, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)* 93+ 29, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*119+169, (2**17)*0+(2**8)*123+ 90, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*132+ 66, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*158+107, (2**17)*0+(2**8)*164+157, (2**17)*0+(2**8)*169+  7, (2**17)*0+(2**8)*181+ 38, (2**17)*0+(2**8)*182+ 48, (2**17)*0+(2**8)*211+ 74, (2**17)*0+(2**8)*231+ 90, (2**17)*0+(2**8)*241+ 81, (2**17)*0+(2**8)*278+155, (2**17)*1+(2**8)*309+ 76, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 12+150, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 31+119, (2**17)*0+(2**8)* 44+150, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 56+ 57, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 76+123, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)* 94+ 49, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*114+  8, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*137+ 28, (2**17)*0+(2**8)*144+ 97, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*150+136, (2**17)*0+(2**8)*165+ 61, (2**17)*0+(2**8)*172+122, (2**17)*0+(2**8)*187+137, (2**17)*0+(2**8)*221+  4, (2**17)*0+(2**8)*249+ 52, (2**17)*0+(2**8)*270+146, (2**17)*1+(2**8)*287+ 63, 
(2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)* 12+ 82, (2**17)*0+(2**8)* 20+154, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 32+149, (2**17)*0+(2**8)* 40+153, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 49+ 64, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*117+121, (2**17)*0+(2**8)*126+  0, (2**17)*0+(2**8)*128+120, (2**17)*0+(2**8)*144+ 36, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*169+ 73, (2**17)*0+(2**8)*179+ 95, (2**17)*0+(2**8)*220+127, (2**17)*0+(2**8)*221+ 33, (2**17)*0+(2**8)*244+156, (2**17)*0+(2**8)*255+  2, (2**17)*0+(2**8)*266+ 31, (2**17)*0+(2**8)*295+133, (2**17)*1+(2**8)*303+156, 
(2**17)*0+(2**8)*  2+ 23, (2**17)*0+(2**8)*  5+ 48, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)*  9+148, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 59+ 88, (2**17)*0+(2**8)* 64+166, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 70+ 25, (2**17)*0+(2**8)* 86+171, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*119+178, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*127+ 85, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*183+151, (2**17)*0+(2**8)*183+ 80, (2**17)*0+(2**8)*214+ 22, (2**17)*0+(2**8)*248+ 53, (2**17)*0+(2**8)*273+143, (2**17)*0+(2**8)*291+166, (2**17)*0+(2**8)*301+165, (2**17)*1+(2**8)*305+ 98, 
(2**17)*0+(2**8)*  0+ 71, (2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 52+163, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 70+123, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*133+127, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*158+143, (2**17)*0+(2**8)*161+134, (2**17)*0+(2**8)*168+ 61, (2**17)*0+(2**8)*189+ 40, (2**17)*0+(2**8)*199+ 99, (2**17)*0+(2**8)*211+ 49, (2**17)*0+(2**8)*220+ 54, (2**17)*0+(2**8)*242+ 76, (2**17)*0+(2**8)*250+160, (2**17)*0+(2**8)*263+ 31, (2**17)*0+(2**8)*267+114, (2**17)*0+(2**8)*290+134, (2**17)*1+(2**8)*311+ 46, 
(2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 13+ 88, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 33+ 49, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 50+ 31, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 80+ 84, (2**17)*0+(2**8)* 88+ 41, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*116+159, (2**17)*0+(2**8)*116+114, (2**17)*0+(2**8)*126+ 83, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*134+ 97, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*166+158, (2**17)*0+(2**8)*174+115, (2**17)*0+(2**8)*193+ 97, (2**17)*0+(2**8)*201+ 48, (2**17)*0+(2**8)*232+ 72, (2**17)*0+(2**8)*238+163, (2**17)*0+(2**8)*308+107, (2**17)*1+(2**8)*315+ 67, 
(2**17)*0+(2**8)*  2+  2, (2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 22+  3, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 42+ 21, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 68+ 98, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 75+110, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)* 93+176, (2**17)*0+(2**8)* 96+ 74, (2**17)*0+(2**8)*100+ 24, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*151+  9, (2**17)*0+(2**8)*154+167, (2**17)*0+(2**8)*167+ 77, (2**17)*0+(2**8)*170+ 49, (2**17)*0+(2**8)*185+ 72, (2**17)*0+(2**8)*209+ 86, (2**17)*0+(2**8)*262+122, (2**17)*0+(2**8)*282+ 68, (2**17)*1+(2**8)*285+  3, 
(2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 11+ 87, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 34+ 89, (2**17)*0+(2**8)* 45+131, (2**17)*0+(2**8)* 48+ 32, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 69+  5, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)* 95+108, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*157+129, (2**17)*0+(2**8)*176+ 30, (2**17)*0+(2**8)*178+170, (2**17)*0+(2**8)*186+ 33, (2**17)*0+(2**8)*222+ 22, (2**17)*0+(2**8)*240+ 76, (2**17)*0+(2**8)*267+173, (2**17)*0+(2**8)*272+137, (2**17)*0+(2**8)*280+ 49, (2**17)*0+(2**8)*299+163, (2**17)*1+(2**8)*302+ 28, 
(2**17)*0+(2**8)*  1+ 87, (2**17)*0+(2**8)*  4+ 29, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 14+ 53, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 32+172, (2**17)*0+(2**8)* 46+  4, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 66+123, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 73+ 40, (2**17)*0+(2**8)* 87+ 48, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)* 97+116, (2**17)*0+(2**8)*100+ 64, (2**17)*0+(2**8)*112+  0, (2**17)*0+(2**8)*118+177, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*133+105, (2**17)*0+(2**8)*150+159, (2**17)*0+(2**8)*152+  0, (2**17)*0+(2**8)*157+149, (2**17)*0+(2**8)*195+116, (2**17)*0+(2**8)*206+ 51, (2**17)*1+(2**8)*299+ 20, 
(2**17)*0+(2**8)*  8+ 15, (2**17)*0+(2**8)* 11+115, (2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 37+ 24, (2**17)*0+(2**8)* 41+ 14, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 54+ 93, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)* 73+ 25, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)* 94+ 90, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*123+ 28, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*147+ 43, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*170+107, (2**17)*0+(2**8)*188+ 63, (2**17)*0+(2**8)*234+ 24, (2**17)*0+(2**8)*247+111, (2**17)*0+(2**8)*263+173, (2**17)*0+(2**8)*272+ 95, (2**17)*0+(2**8)*292+127, (2**17)*1+(2**8)*306+ 72, 
(2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 18+150, (2**17)*0+(2**8)* 31+ 51, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 55+ 34, (2**17)*0+(2**8)* 69+ 77, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 85+ 27, (2**17)*0+(2**8)* 92+ 92, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*124+ 92, (2**17)*0+(2**8)*129+  5, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*140+ 98, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*166+ 93, (2**17)*0+(2**8)*167+179, (2**17)*0+(2**8)*199+ 95, (2**17)*0+(2**8)*202+101, (2**17)*0+(2**8)*224+139, (2**17)*0+(2**8)*270+ 12, (2**17)*0+(2**8)*271+ 54, (2**17)*1+(2**8)*313+ 52, 
(2**17)*0+(2**8)*  6+ 62, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 30+ 13, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 36+ 80, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)* 84+166, (2**17)*0+(2**8)* 85+122, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*147+140, (2**17)*0+(2**8)*152+117, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*160+156, (2**17)*0+(2**8)*174+101, (2**17)*0+(2**8)*207+ 47, (2**17)*0+(2**8)*207+ 62, (2**17)*0+(2**8)*231+ 31, (2**17)*0+(2**8)*235+114, (2**17)*0+(2**8)*266+ 10, (2**17)*0+(2**8)*273+ 40, (2**17)*0+(2**8)*285+ 34, (2**17)*1+(2**8)*298+ 30, 
(2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 53+ 90, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)* 99+143, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*117+ 22, (2**17)*0+(2**8)*126+168, (2**17)*0+(2**8)*129+105, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*159+ 42, (2**17)*0+(2**8)*163+113, (2**17)*0+(2**8)*170+ 43, (2**17)*0+(2**8)*178+165, (2**17)*0+(2**8)*180+129, (2**17)*0+(2**8)*181+109, (2**17)*0+(2**8)*200+ 80, (2**17)*0+(2**8)*227+159, (2**17)*0+(2**8)*227+119, (2**17)*0+(2**8)*256+ 45, (2**17)*0+(2**8)*265+ 73, (2**17)*1+(2**8)*302+165, 
(2**17)*0+(2**8)* 15+168, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 28+165, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 48+ 12, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)* 78+ 60, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)* 98+119, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*124+ 16, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*143+ 36, (2**17)*0+(2**8)*155+ 34, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*162+ 69, (2**17)*0+(2**8)*164+ 81, (2**17)*0+(2**8)*197+ 78, (2**17)*0+(2**8)*217+ 98, (2**17)*0+(2**8)*225+146, (2**17)*0+(2**8)*241+ 89, (2**17)*0+(2**8)*262+115, (2**17)*0+(2**8)*264+ 26, (2**17)*1+(2**8)*281+ 78, 
(2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 19+ 68, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 56+117, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 58+101, (2**17)*0+(2**8)* 68+ 10, (2**17)*0+(2**8)* 77+144, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)* 83+ 81, (2**17)*0+(2**8)* 97+ 80, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*108+115, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*138+  0, (2**17)*0+(2**8)*140+ 69, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*176+150, (2**17)*0+(2**8)*179+148, (2**17)*0+(2**8)*184+168, (2**17)*0+(2**8)*198+155, (2**17)*0+(2**8)*271+139, (2**17)*0+(2**8)*280+159, (2**17)*0+(2**8)*295+ 12, (2**17)*1+(2**8)*301+ 81, 
(2**17)*0+(2**8)*  3+118, (2**17)*0+(2**8)* 11+154, (2**17)*0+(2**8)* 15+ 39, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 52+ 72, (2**17)*0+(2**8)* 58+ 46, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 65+  8, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*130+140, (2**17)*0+(2**8)*138+142, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*159+ 36, (2**17)*0+(2**8)*184+ 19, (2**17)*0+(2**8)*187+ 26, (2**17)*0+(2**8)*222+ 58, (2**17)*0+(2**8)*249+ 53, (2**17)*0+(2**8)*259+ 35, (2**17)*0+(2**8)*261+165, (2**17)*0+(2**8)*264+104, (2**17)*1+(2**8)*306+171, 
(2**17)*0+(2**8)* 17+115, (2**17)*0+(2**8)* 34+ 60, (2**17)*0+(2**8)* 50+ 18, (2**17)*0+(2**8)* 79+ 31, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*161+145, (2**17)*0+(2**8)*175+ 98, (2**17)*0+(2**8)*180+  0, (2**17)*0+(2**8)*185+156, (2**17)*0+(2**8)*200+  0, (2**17)*0+(2**8)*217+119, (2**17)*0+(2**8)*220+  0, (2**17)*0+(2**8)*237+ 15, (2**17)*0+(2**8)*240+  0, (2**17)*0+(2**8)*243+ 11, (2**17)*0+(2**8)*251+168, (2**17)*0+(2**8)*260+  0, (2**17)*0+(2**8)*269+103, (2**17)*0+(2**8)*269+107, (2**17)*0+(2**8)*280+  0, (2**17)*0+(2**8)*281+174, (2**17)*0+(2**8)*296+108, (2**17)*0+(2**8)*300+  0, (2**17)*0+(2**8)*312+ 40, (2**17)*1+(2**8)*313+ 17, 
(2**17)*0+(2**8)* 17+ 59, (2**17)*0+(2**8)* 35+ 24, (2**17)*0+(2**8)* 59+153, (2**17)*0+(2**8)* 63+ 26, (2**17)*0+(2**8)* 66+145, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*163+174, (2**17)*0+(2**8)*168+ 94, (2**17)*0+(2**8)*181+  0, (2**17)*0+(2**8)*190+164, (2**17)*0+(2**8)*201+  0, (2**17)*0+(2**8)*203+ 40, (2**17)*0+(2**8)*221+  0, (2**17)*0+(2**8)*241+  0, (2**17)*0+(2**8)*246+ 37, (2**17)*0+(2**8)*252+113, (2**17)*0+(2**8)*261+  0, (2**17)*0+(2**8)*268+ 56, (2**17)*0+(2**8)*275+165, (2**17)*0+(2**8)*281+  0, (2**17)*0+(2**8)*296+153, (2**17)*0+(2**8)*297+ 99, (2**17)*0+(2**8)*301+  0, (2**17)*0+(2**8)*314+ 45, (2**17)*1+(2**8)*316+ 42, 
(2**17)*0+(2**8)*  0+ 80, (2**17)*0+(2**8)*  7+158, (2**17)*0+(2**8)* 29+130, (2**17)*0+(2**8)* 43+140, (2**17)*0+(2**8)* 55+117, (2**17)*0+(2**8)* 72+174, (2**17)*0+(2**8)* 91+ 90, (2**17)*0+(2**8)*101+ 51, (2**17)*0+(2**8)*122+176, (2**17)*0+(2**8)*128+ 61, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*177+ 37, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*198+ 95, (2**17)*0+(2**8)*202+  0, (2**17)*0+(2**8)*222+  0, (2**17)*0+(2**8)*236+121, (2**17)*0+(2**8)*242+  0, (2**17)*0+(2**8)*258+ 44, (2**17)*0+(2**8)*262+  0, (2**17)*0+(2**8)*265+ 59, (2**17)*0+(2**8)*282+  0, (2**17)*0+(2**8)*302+  0, (2**17)*0+(2**8)*308+130, (2**17)*1+(2**8)*309+118, 
(2**17)*0+(2**8)* 13+ 33, (2**17)*0+(2**8)* 26+ 58, (2**17)*0+(2**8)* 45+144, (2**17)*0+(2**8)* 63+ 86, (2**17)*0+(2**8)* 79+122, (2**17)*0+(2**8)* 82+ 14, (2**17)*0+(2**8)*115+129, (2**17)*0+(2**8)*134+ 86, (2**17)*0+(2**8)*156+ 61, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*165+ 92, (2**17)*0+(2**8)*173+148, (2**17)*0+(2**8)*183+  0, (2**17)*0+(2**8)*196+104, (2**17)*0+(2**8)*203+  0, (2**17)*0+(2**8)*213+ 56, (2**17)*0+(2**8)*223+  0, (2**17)*0+(2**8)*243+  0, (2**17)*0+(2**8)*250+100, (2**17)*0+(2**8)*263+  0, (2**17)*0+(2**8)*274+ 35, (2**17)*0+(2**8)*283+  0, (2**17)*0+(2**8)*291+156, (2**17)*0+(2**8)*303+  0, (2**17)*1+(2**8)*305+101, 
(2**17)*0+(2**8)*  4+156, (2**17)*0+(2**8)*  9+  6, (2**17)*0+(2**8)* 21+ 37, (2**17)*0+(2**8)* 22+ 47, (2**17)*0+(2**8)* 51+ 73, (2**17)*0+(2**8)* 71+ 89, (2**17)*0+(2**8)* 81+ 80, (2**17)*0+(2**8)*118+154, (2**17)*0+(2**8)*149+ 75, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*176+ 41, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*204+  0, (2**17)*0+(2**8)*204+ 13, (2**17)*0+(2**8)*224+  0, (2**17)*0+(2**8)*234+124, (2**17)*0+(2**8)*244+  0, (2**17)*0+(2**8)*253+ 29, (2**17)*0+(2**8)*264+  0, (2**17)*0+(2**8)*279+169, (2**17)*0+(2**8)*283+ 90, (2**17)*0+(2**8)*284+  0, (2**17)*0+(2**8)*292+ 66, (2**17)*0+(2**8)*304+  0, (2**17)*1+(2**8)*318+107, 
(2**17)*0+(2**8)*  5+ 60, (2**17)*0+(2**8)* 12+121, (2**17)*0+(2**8)* 27+136, (2**17)*0+(2**8)* 61+  3, (2**17)*0+(2**8)* 89+ 51, (2**17)*0+(2**8)*110+145, (2**17)*0+(2**8)*127+ 62, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*172+150, (2**17)*0+(2**8)*185+  0, (2**17)*0+(2**8)*191+119, (2**17)*0+(2**8)*204+150, (2**17)*0+(2**8)*205+  0, (2**17)*0+(2**8)*216+ 57, (2**17)*0+(2**8)*225+  0, (2**17)*0+(2**8)*236+123, (2**17)*0+(2**8)*245+  0, (2**17)*0+(2**8)*254+ 49, (2**17)*0+(2**8)*265+  0, (2**17)*0+(2**8)*274+  8, (2**17)*0+(2**8)*285+  0, (2**17)*0+(2**8)*297+ 28, (2**17)*0+(2**8)*304+ 97, (2**17)*0+(2**8)*305+  0, (2**17)*1+(2**8)*310+136, 
(2**17)*0+(2**8)*  9+ 72, (2**17)*0+(2**8)* 19+ 94, (2**17)*0+(2**8)* 60+126, (2**17)*0+(2**8)* 61+ 32, (2**17)*0+(2**8)* 84+155, (2**17)*0+(2**8)* 95+  1, (2**17)*0+(2**8)*106+ 30, (2**17)*0+(2**8)*135+132, (2**17)*0+(2**8)*143+155, (2**17)*0+(2**8)*166+  0, (2**17)*0+(2**8)*172+ 82, (2**17)*0+(2**8)*180+154, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*192+149, (2**17)*0+(2**8)*200+153, (2**17)*0+(2**8)*206+  0, (2**17)*0+(2**8)*209+ 64, (2**17)*0+(2**8)*226+  0, (2**17)*0+(2**8)*246+  0, (2**17)*0+(2**8)*266+  0, (2**17)*0+(2**8)*277+121, (2**17)*0+(2**8)*286+  0, (2**17)*0+(2**8)*288+120, (2**17)*0+(2**8)*304+ 36, (2**17)*1+(2**8)*306+  0, 
(2**17)*0+(2**8)* 23+150, (2**17)*0+(2**8)* 23+ 79, (2**17)*0+(2**8)* 54+ 21, (2**17)*0+(2**8)* 88+ 52, (2**17)*0+(2**8)*113+142, (2**17)*0+(2**8)*131+165, (2**17)*0+(2**8)*141+164, (2**17)*0+(2**8)*145+ 97, (2**17)*0+(2**8)*162+ 23, (2**17)*0+(2**8)*165+ 48, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*169+148, (2**17)*0+(2**8)*187+  0, (2**17)*0+(2**8)*207+  0, (2**17)*0+(2**8)*219+ 88, (2**17)*0+(2**8)*224+166, (2**17)*0+(2**8)*227+  0, (2**17)*0+(2**8)*230+ 25, (2**17)*0+(2**8)*246+171, (2**17)*0+(2**8)*247+  0, (2**17)*0+(2**8)*267+  0, (2**17)*0+(2**8)*279+178, (2**17)*0+(2**8)*287+  0, (2**17)*0+(2**8)*287+ 85, (2**17)*1+(2**8)*307+  0, 
(2**17)*0+(2**8)*  1+133, (2**17)*0+(2**8)*  8+ 60, (2**17)*0+(2**8)* 29+ 39, (2**17)*0+(2**8)* 39+ 98, (2**17)*0+(2**8)* 51+ 48, (2**17)*0+(2**8)* 60+ 53, (2**17)*0+(2**8)* 82+ 75, (2**17)*0+(2**8)* 90+159, (2**17)*0+(2**8)*103+ 30, (2**17)*0+(2**8)*107+113, (2**17)*0+(2**8)*130+133, (2**17)*0+(2**8)*151+ 45, (2**17)*0+(2**8)*160+ 71, (2**17)*0+(2**8)*168+  0, (2**17)*0+(2**8)*188+  0, (2**17)*0+(2**8)*208+  0, (2**17)*0+(2**8)*212+163, (2**17)*0+(2**8)*228+  0, (2**17)*0+(2**8)*230+123, (2**17)*0+(2**8)*248+  0, (2**17)*0+(2**8)*268+  0, (2**17)*0+(2**8)*288+  0, (2**17)*0+(2**8)*293+127, (2**17)*0+(2**8)*308+  0, (2**17)*1+(2**8)*318+143, 
(2**17)*0+(2**8)*  6+157, (2**17)*0+(2**8)* 14+114, (2**17)*0+(2**8)* 33+ 96, (2**17)*0+(2**8)* 41+ 47, (2**17)*0+(2**8)* 72+ 71, (2**17)*0+(2**8)* 78+162, (2**17)*0+(2**8)*148+106, (2**17)*0+(2**8)*155+ 66, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*173+ 88, (2**17)*0+(2**8)*189+  0, (2**17)*0+(2**8)*193+ 49, (2**17)*0+(2**8)*209+  0, (2**17)*0+(2**8)*210+ 31, (2**17)*0+(2**8)*229+  0, (2**17)*0+(2**8)*240+ 84, (2**17)*0+(2**8)*248+ 41, (2**17)*0+(2**8)*249+  0, (2**17)*0+(2**8)*269+  0, (2**17)*0+(2**8)*276+159, (2**17)*0+(2**8)*276+114, (2**17)*0+(2**8)*286+ 83, (2**17)*0+(2**8)*289+  0, (2**17)*0+(2**8)*294+ 97, (2**17)*1+(2**8)*309+  0, 
(2**17)*0+(2**8)*  7+ 76, (2**17)*0+(2**8)* 10+ 48, (2**17)*0+(2**8)* 25+ 71, (2**17)*0+(2**8)* 49+ 85, (2**17)*0+(2**8)*102+121, (2**17)*0+(2**8)*122+ 67, (2**17)*0+(2**8)*125+  2, (2**17)*0+(2**8)*162+  2, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*182+  3, (2**17)*0+(2**8)*190+  0, (2**17)*0+(2**8)*202+ 21, (2**17)*0+(2**8)*210+  0, (2**17)*0+(2**8)*228+ 98, (2**17)*0+(2**8)*230+  0, (2**17)*0+(2**8)*235+110, (2**17)*0+(2**8)*250+  0, (2**17)*0+(2**8)*253+176, (2**17)*0+(2**8)*256+ 74, (2**17)*0+(2**8)*260+ 24, (2**17)*0+(2**8)*270+  0, (2**17)*0+(2**8)*290+  0, (2**17)*0+(2**8)*310+  0, (2**17)*0+(2**8)*311+  9, (2**17)*1+(2**8)*314+167, 
(2**17)*0+(2**8)* 16+ 29, (2**17)*0+(2**8)* 18+169, (2**17)*0+(2**8)* 26+ 32, (2**17)*0+(2**8)* 62+ 21, (2**17)*0+(2**8)* 80+ 75, (2**17)*0+(2**8)*107+172, (2**17)*0+(2**8)*112+136, (2**17)*0+(2**8)*120+ 48, (2**17)*0+(2**8)*139+162, (2**17)*0+(2**8)*142+ 27, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*171+ 87, (2**17)*0+(2**8)*191+  0, (2**17)*0+(2**8)*194+ 89, (2**17)*0+(2**8)*205+131, (2**17)*0+(2**8)*208+ 32, (2**17)*0+(2**8)*211+  0, (2**17)*0+(2**8)*229+  5, (2**17)*0+(2**8)*231+  0, (2**17)*0+(2**8)*251+  0, (2**17)*0+(2**8)*255+108, (2**17)*0+(2**8)*271+  0, (2**17)*0+(2**8)*291+  0, (2**17)*0+(2**8)*311+  0, (2**17)*1+(2**8)*317+129, 
(2**17)*0+(2**8)* 35+115, (2**17)*0+(2**8)* 46+ 50, (2**17)*0+(2**8)*139+ 19, (2**17)*0+(2**8)*161+ 87, (2**17)*0+(2**8)*164+ 29, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*174+ 53, (2**17)*0+(2**8)*192+  0, (2**17)*0+(2**8)*192+172, (2**17)*0+(2**8)*206+  4, (2**17)*0+(2**8)*212+  0, (2**17)*0+(2**8)*226+123, (2**17)*0+(2**8)*232+  0, (2**17)*0+(2**8)*233+ 40, (2**17)*0+(2**8)*247+ 48, (2**17)*0+(2**8)*252+  0, (2**17)*0+(2**8)*257+116, (2**17)*0+(2**8)*260+ 64, (2**17)*0+(2**8)*272+  0, (2**17)*0+(2**8)*278+177, (2**17)*0+(2**8)*292+  0, (2**17)*0+(2**8)*293+105, (2**17)*0+(2**8)*310+159, (2**17)*0+(2**8)*312+  0, (2**17)*1+(2**8)*317+149, 
(2**17)*0+(2**8)* 10+106, (2**17)*0+(2**8)* 28+ 62, (2**17)*0+(2**8)* 74+ 23, (2**17)*0+(2**8)* 87+110, (2**17)*0+(2**8)*103+172, (2**17)*0+(2**8)*112+ 94, (2**17)*0+(2**8)*132+126, (2**17)*0+(2**8)*146+ 71, (2**17)*0+(2**8)*168+ 15, (2**17)*0+(2**8)*171+115, (2**17)*0+(2**8)*173+  0, (2**17)*0+(2**8)*193+  0, (2**17)*0+(2**8)*197+ 24, (2**17)*0+(2**8)*201+ 14, (2**17)*0+(2**8)*213+  0, (2**17)*0+(2**8)*214+ 93, (2**17)*0+(2**8)*233+  0, (2**17)*0+(2**8)*233+ 25, (2**17)*0+(2**8)*253+  0, (2**17)*0+(2**8)*254+ 90, (2**17)*0+(2**8)*273+  0, (2**17)*0+(2**8)*283+ 28, (2**17)*0+(2**8)*293+  0, (2**17)*0+(2**8)*307+ 43, (2**17)*1+(2**8)*313+  0, 
(2**17)*0+(2**8)*  6+ 92, (2**17)*0+(2**8)*  7+178, (2**17)*0+(2**8)* 39+ 94, (2**17)*0+(2**8)* 42+100, (2**17)*0+(2**8)* 64+138, (2**17)*0+(2**8)*110+ 11, (2**17)*0+(2**8)*111+ 53, (2**17)*0+(2**8)*153+ 51, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*178+150, (2**17)*0+(2**8)*191+ 51, (2**17)*0+(2**8)*194+  0, (2**17)*0+(2**8)*214+  0, (2**17)*0+(2**8)*215+ 34, (2**17)*0+(2**8)*229+ 77, (2**17)*0+(2**8)*234+  0, (2**17)*0+(2**8)*245+ 27, (2**17)*0+(2**8)*252+ 92, (2**17)*0+(2**8)*254+  0, (2**17)*0+(2**8)*274+  0, (2**17)*0+(2**8)*284+ 92, (2**17)*0+(2**8)*289+  5, (2**17)*0+(2**8)*294+  0, (2**17)*0+(2**8)*300+ 98, (2**17)*1+(2**8)*314+  0, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)* 14+100, (2**17)*0+(2**8)* 47+ 46, (2**17)*0+(2**8)* 47+ 61, (2**17)*0+(2**8)* 71+ 30, (2**17)*0+(2**8)* 75+113, (2**17)*0+(2**8)*106+  9, (2**17)*0+(2**8)*113+ 39, (2**17)*0+(2**8)*125+ 33, (2**17)*0+(2**8)*138+ 29, (2**17)*0+(2**8)*166+ 62, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*190+ 13, (2**17)*0+(2**8)*195+  0, (2**17)*0+(2**8)*196+ 80, (2**17)*0+(2**8)*215+  0, (2**17)*0+(2**8)*235+  0, (2**17)*0+(2**8)*244+166, (2**17)*0+(2**8)*245+122, (2**17)*0+(2**8)*255+  0, (2**17)*0+(2**8)*275+  0, (2**17)*0+(2**8)*295+  0, (2**17)*0+(2**8)*307+140, (2**17)*0+(2**8)*312+117, (2**17)*1+(2**8)*315+  0, 
(2**17)*0+(2**8)*  3+112, (2**17)*0+(2**8)* 10+ 42, (2**17)*0+(2**8)* 18+164, (2**17)*0+(2**8)* 20+128, (2**17)*0+(2**8)* 21+108, (2**17)*0+(2**8)* 40+ 79, (2**17)*0+(2**8)* 67+158, (2**17)*0+(2**8)* 67+118, (2**17)*0+(2**8)* 96+ 44, (2**17)*0+(2**8)*105+ 72, (2**17)*0+(2**8)*142+164, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*213+ 90, (2**17)*0+(2**8)*216+  0, (2**17)*0+(2**8)*236+  0, (2**17)*0+(2**8)*256+  0, (2**17)*0+(2**8)*259+143, (2**17)*0+(2**8)*276+  0, (2**17)*0+(2**8)*277+ 22, (2**17)*0+(2**8)*286+168, (2**17)*0+(2**8)*289+105, (2**17)*0+(2**8)*296+  0, (2**17)*0+(2**8)*316+  0, (2**17)*1+(2**8)*319+ 42, 
(2**17)*0+(2**8)*  2+ 68, (2**17)*0+(2**8)*  4+ 80, (2**17)*0+(2**8)* 37+ 77, (2**17)*0+(2**8)* 57+ 97, (2**17)*0+(2**8)* 65+145, (2**17)*0+(2**8)* 81+ 88, (2**17)*0+(2**8)*102+114, (2**17)*0+(2**8)*104+ 25, (2**17)*0+(2**8)*121+ 77, (2**17)*0+(2**8)*175+168, (2**17)*0+(2**8)*177+  0, (2**17)*0+(2**8)*188+165, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*208+ 12, (2**17)*0+(2**8)*217+  0, (2**17)*0+(2**8)*237+  0, (2**17)*0+(2**8)*238+ 60, (2**17)*0+(2**8)*257+  0, (2**17)*0+(2**8)*258+119, (2**17)*0+(2**8)*277+  0, (2**17)*0+(2**8)*284+ 16, (2**17)*0+(2**8)*297+  0, (2**17)*0+(2**8)*303+ 36, (2**17)*0+(2**8)*315+ 34, (2**17)*1+(2**8)*317+  0, 
(2**17)*0+(2**8)* 16+149, (2**17)*0+(2**8)* 19+147, (2**17)*0+(2**8)* 24+167, (2**17)*0+(2**8)* 38+154, (2**17)*0+(2**8)*111+138, (2**17)*0+(2**8)*120+158, (2**17)*0+(2**8)*135+ 11, (2**17)*0+(2**8)*141+ 80, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*179+ 68, (2**17)*0+(2**8)*198+  0, (2**17)*0+(2**8)*216+117, (2**17)*0+(2**8)*218+  0, (2**17)*0+(2**8)*218+101, (2**17)*0+(2**8)*228+ 10, (2**17)*0+(2**8)*237+144, (2**17)*0+(2**8)*238+  0, (2**17)*0+(2**8)*243+ 81, (2**17)*0+(2**8)*257+ 80, (2**17)*0+(2**8)*258+  0, (2**17)*0+(2**8)*268+115, (2**17)*0+(2**8)*278+  0, (2**17)*0+(2**8)*298+  0, (2**17)*0+(2**8)*300+ 69, (2**17)*1+(2**8)*318+  0, 
(2**17)*0+(2**8)* 24+ 18, (2**17)*0+(2**8)* 27+ 25, (2**17)*0+(2**8)* 62+ 57, (2**17)*0+(2**8)* 89+ 52, (2**17)*0+(2**8)* 99+ 34, (2**17)*0+(2**8)*101+164, (2**17)*0+(2**8)*104+103, (2**17)*0+(2**8)*146+170, (2**17)*0+(2**8)*163+118, (2**17)*0+(2**8)*171+154, (2**17)*0+(2**8)*175+ 39, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*199+  0, (2**17)*0+(2**8)*212+ 72, (2**17)*0+(2**8)*218+ 46, (2**17)*0+(2**8)*219+  0, (2**17)*0+(2**8)*225+  8, (2**17)*0+(2**8)*239+  0, (2**17)*0+(2**8)*259+  0, (2**17)*0+(2**8)*279+  0, (2**17)*0+(2**8)*290+140, (2**17)*0+(2**8)*298+142, (2**17)*0+(2**8)*299+  0, (2**17)*0+(2**8)*319+  0, (2**17)*1+(2**8)*319+ 36, 


(2**17)*0+(2**8)*  0+  0, (2**17)*0+(2**8)*  1+145, (2**17)*0+(2**8)* 11+150, (2**17)*0+(2**8)* 13+ 98, (2**17)*0+(2**8)* 18+  0, (2**17)*0+(2**8)* 26+156, (2**17)*0+(2**8)* 36+  0, (2**17)*0+(2**8)* 37+104, (2**17)*0+(2**8)* 53+ 63, (2**17)*0+(2**8)* 54+  0, (2**17)*0+(2**8)* 57+ 57, (2**17)*0+(2**8)* 72+  0, (2**17)*0+(2**8)* 84+ 37, (2**17)*0+(2**8)* 90+  0, (2**17)*0+(2**8)* 91+  4, (2**17)*0+(2**8)*108+  0, (2**17)*0+(2**8)*112+174, (2**17)*0+(2**8)*124+108, (2**17)*0+(2**8)*126+  0, (2**17)*0+(2**8)*126+ 47, (2**17)*0+(2**8)*131+ 29, (2**17)*0+(2**8)*144+  0, (2**17)*0+(2**8)*154+ 32, (2**17)*0+(2**8)*197+ 61, (2**17)*0+(2**8)*226+146, (2**17)*0+(2**8)*248+ 52, (2**17)*0+(2**8)*259+119, (2**17)*1+(2**8)*315+ 33, 
(2**17)*0+(2**8)*  1+  0, (2**17)*0+(2**8)*  3+174, (2**17)*0+(2**8)*  7+ 94, (2**17)*0+(2**8)* 12+148, (2**17)*0+(2**8)* 19+  0, (2**17)*0+(2**8)* 31+164, (2**17)*0+(2**8)* 37+  0, (2**17)*0+(2**8)* 44+ 40, (2**17)*0+(2**8)* 55+  0, (2**17)*0+(2**8)* 73+  0, (2**17)*0+(2**8)* 75+ 15, (2**17)*0+(2**8)* 87+100, (2**17)*0+(2**8)* 91+  0, (2**17)*0+(2**8)*100+107, (2**17)*0+(2**8)*109+  0, (2**17)*0+(2**8)*118+148, (2**17)*0+(2**8)*119+ 18, (2**17)*0+(2**8)*127+  0, (2**17)*0+(2**8)*140+ 18, (2**17)*0+(2**8)*143+117, (2**17)*0+(2**8)*145+  0, (2**17)*0+(2**8)*158+150, (2**17)*0+(2**8)*192+131, (2**17)*0+(2**8)*206+141, (2**17)*0+(2**8)*218+118, (2**17)*0+(2**8)*224+ 87, (2**17)*0+(2**8)*256+ 52, (2**17)*1+(2**8)*306+161, 
(2**17)*0+(2**8)*  2+  0, (2**17)*0+(2**8)* 16+ 37, (2**17)*0+(2**8)* 20+  0, (2**17)*0+(2**8)* 38+  0, (2**17)*0+(2**8)* 56+  0, (2**17)*0+(2**8)* 58+119, (2**17)*0+(2**8)* 74+  0, (2**17)*0+(2**8)* 92+  0, (2**17)*0+(2**8)* 98+ 56, (2**17)*0+(2**8)*100+103, (2**17)*0+(2**8)*110+  0, (2**17)*0+(2**8)*124+153, (2**17)*0+(2**8)*128+  0, (2**17)*0+(2**8)*137+130, (2**17)*0+(2**8)*143+ 40, (2**17)*0+(2**8)*146+  0, (2**17)*0+(2**8)*146+ 42, (2**17)*0+(2**8)*159+141, (2**17)*0+(2**8)*162+ 81, (2**17)*0+(2**8)*170+  7, (2**17)*0+(2**8)*189+ 59, (2**17)*0+(2**8)*196+ 97, (2**17)*0+(2**8)*198+ 25, (2**17)*0+(2**8)*202+ 95, (2**17)*0+(2**8)*224+ 27, (2**17)*0+(2**8)*241+115, (2**17)*0+(2**8)*244+122, (2**17)*1+(2**8)*271+145, 
(2**17)*0+(2**8)*  3+  0, (2**17)*0+(2**8)*  5+ 92, (2**17)*0+(2**8)* 21+  0, (2**17)*0+(2**8)* 39+  0, (2**17)*0+(2**8)* 39+ 95, (2**17)*0+(2**8)* 57+  0, (2**17)*0+(2**8)* 71+ 25, (2**17)*0+(2**8)* 75+  0, (2**17)*0+(2**8)* 79+ 30, (2**17)*0+(2**8)* 93+  0, (2**17)*0+(2**8)*105+ 35, (2**17)*0+(2**8)*108+ 88, (2**17)*0+(2**8)*111+  0, (2**17)*0+(2**8)*129+  0, (2**17)*0+(2**8)*135+101, (2**17)*0+(2**8)*147+  0, (2**17)*0+(2**8)*174+ 34, (2**17)*0+(2**8)*178+ 60, (2**17)*0+(2**8)*182+ 95, (2**17)*0+(2**8)*185+ 48, (2**17)*0+(2**8)*214+ 19, (2**17)*0+(2**8)*231+ 90, (2**17)*0+(2**8)*240+ 15, (2**17)*0+(2**8)*268+130, (2**17)*0+(2**8)*272+155, (2**17)*0+(2**8)*300+ 85, (2**17)*0+(2**8)*308+ 62, (2**17)*1+(2**8)*314+ 38, 
(2**17)*0+(2**8)*  4+  0, (2**17)*0+(2**8)* 14+ 41, (2**17)*0+(2**8)* 22+  0, (2**17)*0+(2**8)* 40+  0, (2**17)*0+(2**8)* 51+ 64, (2**17)*0+(2**8)* 58+  0, (2**17)*0+(2**8)* 68+123, (2**17)*0+(2**8)* 76+  0, (2**17)*0+(2**8)* 90+ 49, (2**17)*0+(2**8)* 90+ 90, (2**17)*0+(2**8)* 94+  0, (2**17)*0+(2**8)*112+  0, (2**17)*0+(2**8)*114+ 90, (2**17)*0+(2**8)*126+162, (2**17)*0+(2**8)*130+  0, (2**17)*0+(2**8)*134+ 97, (2**17)*0+(2**8)*148+  0, (2**17)*0+(2**8)*155+149, (2**17)*0+(2**8)*166+157, (2**17)*0+(2**8)*167+ 61, (2**17)*0+(2**8)*184+ 38, (2**17)*0+(2**8)*186+ 80, (2**17)*0+(2**8)*207+ 17, (2**17)*0+(2**8)*223+ 33, (2**17)*0+(2**8)*239+ 81, (2**17)*0+(2**8)*242+ 65, (2**17)*0+(2**8)*277+112, (2**17)*1+(2**8)*314+139, 
(2**17)*0+(2**8)*  5+  0, (2**17)*0+(2**8)* 11+ 82, (2**17)*0+(2**8)* 18+150, (2**17)*0+(2**8)* 23+  0, (2**17)*0+(2**8)* 32+119, (2**17)*0+(2**8)* 41+  0, (2**17)*0+(2**8)* 46+150, (2**17)*0+(2**8)* 46+ 13, (2**17)*0+(2**8)* 59+  0, (2**17)*0+(2**8)* 74+123, (2**17)*0+(2**8)* 74+121, (2**17)*0+(2**8)* 77+  0, (2**17)*0+(2**8)* 92+ 44, (2**17)*0+(2**8)* 95+  0, (2**17)*0+(2**8)*105+  8, (2**17)*0+(2**8)*113+  0, (2**17)*0+(2**8)*131+  0, (2**17)*0+(2**8)*149+  0, (2**17)*0+(2**8)*149+ 42, (2**17)*0+(2**8)*170+ 73, (2**17)*0+(2**8)*178+116, (2**17)*0+(2**8)*221+154, (2**17)*0+(2**8)*223+  4, (2**17)*0+(2**8)*283+106, (2**17)*0+(2**8)*284+ 87, (2**17)*0+(2**8)*294+176, (2**17)*0+(2**8)*295+156, (2**17)*1+(2**8)*321+ 75, 
(2**17)*0+(2**8)*  2+ 23, (2**17)*0+(2**8)*  5+ 48, (2**17)*0+(2**8)*  6+  0, (2**17)*0+(2**8)*  8+148, (2**17)*0+(2**8)* 19+ 83, (2**17)*0+(2**8)* 21+154, (2**17)*0+(2**8)* 24+  0, (2**17)*0+(2**8)* 42+  0, (2**17)*0+(2**8)* 52+ 31, (2**17)*0+(2**8)* 60+  0, (2**17)*0+(2**8)* 68+ 25, (2**17)*0+(2**8)* 78+  0, (2**17)*0+(2**8)* 93+143, (2**17)*0+(2**8)* 95+ 75, (2**17)*0+(2**8)* 96+  0, (2**17)*0+(2**8)*114+  0, (2**17)*0+(2**8)*132+  0, (2**17)*0+(2**8)*148+107, (2**17)*0+(2**8)*150+  0, (2**17)*0+(2**8)*202+ 99, (2**17)*0+(2**8)*222+127, (2**17)*0+(2**8)*240+ 76, (2**17)*0+(2**8)*249+160, (2**17)*0+(2**8)*275+ 73, (2**17)*0+(2**8)*283+140, (2**17)*0+(2**8)*297+ 98, (2**17)*0+(2**8)*301+ 73, (2**17)*1+(2**8)*313+147, 
(2**17)*0+(2**8)*  0+ 71, (2**17)*0+(2**8)*  7+  0, (2**17)*0+(2**8)* 25+  0, (2**17)*0+(2**8)* 41+153, (2**17)*0+(2**8)* 43+  0, (2**17)*0+(2**8)* 56+ 34, (2**17)*0+(2**8)* 61+  0, (2**17)*0+(2**8)* 79+  0, (2**17)*0+(2**8)* 84+171, (2**17)*0+(2**8)* 92+119, (2**17)*0+(2**8)* 97+  0, (2**17)*0+(2**8)*115+  0, (2**17)*0+(2**8)*116+ 85, (2**17)*0+(2**8)*133+  0, (2**17)*0+(2**8)*134+ 36, (2**17)*0+(2**8)*148+143, (2**17)*0+(2**8)*151+  0, (2**17)*0+(2**8)*156+ 39, (2**17)*0+(2**8)*163+134, (2**17)*0+(2**8)*169+ 61, (2**17)*0+(2**8)*186+151, (2**17)*0+(2**8)*190+137, (2**17)*0+(2**8)*198+116, (2**17)*0+(2**8)*220+ 98, (2**17)*0+(2**8)*243+156, (2**17)*0+(2**8)*253+ 60, (2**17)*0+(2**8)*278+ 63, (2**17)*1+(2**8)*298+ 64, 
(2**17)*0+(2**8)*  8+  0, (2**17)*0+(2**8)* 17+  7, (2**17)*0+(2**8)* 26+  0, (2**17)*0+(2**8)* 44+  0, (2**17)*0+(2**8)* 47+131, (2**17)*0+(2**8)* 62+  0, (2**17)*0+(2**8)* 63+ 30, (2**17)*0+(2**8)* 80+  0, (2**17)*0+(2**8)* 88+168, (2**17)*0+(2**8)* 98+  0, (2**17)*0+(2**8)*107+177, (2**17)*0+(2**8)*116+  0, (2**17)*0+(2**8)*118+ 33, (2**17)*0+(2**8)*131+ 41, (2**17)*0+(2**8)*134+  0, (2**17)*0+(2**8)*141+173, (2**17)*0+(2**8)*152+  0, (2**17)*0+(2**8)*161+ 94, (2**17)*0+(2**8)*168+158, (2**17)*0+(2**8)*173+122, (2**17)*0+(2**8)*188+ 72, (2**17)*0+(2**8)*192+ 40, (2**17)*0+(2**8)*209+145, (2**17)*0+(2**8)*217+ 22, (2**17)*0+(2**8)*250+ 91, (2**17)*0+(2**8)*264+171, (2**17)*0+(2**8)*271+ 59, (2**17)*1+(2**8)*312+ 88, 
(2**17)*0+(2**8)*  2+  2, (2**17)*0+(2**8)*  9+  0, (2**17)*0+(2**8)* 23+  3, (2**17)*0+(2**8)* 27+  0, (2**17)*0+(2**8)* 43+ 21, (2**17)*0+(2**8)* 45+  0, (2**17)*0+(2**8)* 63+  0, (2**17)*0+(2**8)* 81+  0, (2**17)*0+(2**8)* 97+ 19, (2**17)*0+(2**8)* 99+  0, (2**17)*0+(2**8)*106+165, (2**17)*0+(2**8)*117+  0, (2**17)*0+(2**8)*120+127, (2**17)*0+(2**8)*128+171, (2**17)*0+(2**8)*135+  0, (2**17)*0+(2**8)*153+  0, (2**17)*0+(2**8)*171+ 49, (2**17)*0+(2**8)*177+107, (2**17)*0+(2**8)*189+ 33, (2**17)*0+(2**8)*204+ 48, (2**17)*0+(2**8)*222+ 54, (2**17)*0+(2**8)*232+ 72, (2**17)*0+(2**8)*234+ 24, (2**17)*0+(2**8)*242+167, (2**17)*0+(2**8)*285+133, (2**17)*0+(2**8)*302+ 91, (2**17)*0+(2**8)*307+ 67, (2**17)*1+(2**8)*322+ 49, 
(2**17)*0+(2**8)* 10+  0, (2**17)*0+(2**8)* 10+ 87, (2**17)*0+(2**8)* 28+  0, (2**17)*0+(2**8)* 32+ 51, (2**17)*0+(2**8)* 33+149, (2**17)*0+(2**8)* 38+ 24, (2**17)*0+(2**8)* 46+  0, (2**17)*0+(2**8)* 54+163, (2**17)*0+(2**8)* 64+  0, (2**17)*0+(2**8)* 67+ 77, (2**17)*0+(2**8)* 73+110, (2**17)*0+(2**8)* 82+  0, (2**17)*0+(2**8)* 89+ 92, (2**17)*0+(2**8)*100+  0, (2**17)*0+(2**8)*108+130, (2**17)*0+(2**8)*114+ 28, (2**17)*0+(2**8)*118+  0, (2**17)*0+(2**8)*132+112, (2**17)*0+(2**8)*136+  0, (2**17)*0+(2**8)*139+ 78, (2**17)*0+(2**8)*154+  0, (2**17)*0+(2**8)*154+121, (2**17)*0+(2**8)*176+ 30, (2**17)*0+(2**8)*179+ 66, (2**17)*0+(2**8)*213+ 86, (2**17)*0+(2**8)*255+ 35, (2**17)*0+(2**8)*266+143, (2**17)*1+(2**8)*322+  9, 
(2**17)*0+(2**8)*  1+ 87, (2**17)*0+(2**8)*  4+ 29, (2**17)*0+(2**8)* 11+  0, (2**17)*0+(2**8)* 12+ 88, (2**17)*0+(2**8)* 29+  0, (2**17)*0+(2**8)* 34+ 49, (2**17)*0+(2**8)* 47+  0, (2**17)*0+(2**8)* 48+  4, (2**17)*0+(2**8)* 55+ 93, (2**17)*0+(2**8)* 65+  0, (2**17)*0+(2**8)* 67+  5, (2**17)*0+(2**8)* 72+124, (2**17)*0+(2**8)* 83+  0, (2**17)*0+(2**8)*101+  0, (2**17)*0+(2**8)*101+142, (2**17)*0+(2**8)*102+ 92, (2**17)*0+(2**8)*119+  0, (2**17)*0+(2**8)*120+105, (2**17)*0+(2**8)*137+  0, (2**17)*0+(2**8)*155+  0, (2**17)*0+(2**8)*161+ 55, (2**17)*0+(2**8)*191+ 63, (2**17)*0+(2**8)*200+ 78, (2**17)*0+(2**8)*235+114, (2**17)*0+(2**8)*273+ 49, (2**17)*0+(2**8)*292+ 62, (2**17)*0+(2**8)*299+107, (2**17)*1+(2**8)*309+156, 
(2**17)*0+(2**8)*  7+ 15, (2**17)*0+(2**8)* 12+  0, (2**17)*0+(2**8)* 30+  0, (2**17)*0+(2**8)* 31+ 13, (2**17)*0+(2**8)* 35+ 89, (2**17)*0+(2**8)* 42+ 14, (2**17)*0+(2**8)* 48+  0, (2**17)*0+(2**8)* 50+ 32, (2**17)*0+(2**8)* 64+123, (2**17)*0+(2**8)* 66+  0, (2**17)*0+(2**8)* 66+ 98, (2**17)*0+(2**8)* 83+ 27, (2**17)*0+(2**8)* 84+  0, (2**17)*0+(2**8)* 96+ 93, (2**17)*0+(2**8)*102+  0, (2**17)*0+(2**8)*107+126, (2**17)*0+(2**8)*110+177, (2**17)*0+(2**8)*120+  0, (2**17)*0+(2**8)*129+ 98, (2**17)*0+(2**8)*130+176, (2**17)*0+(2**8)*138+  0, (2**17)*0+(2**8)*144+ 44, (2**17)*0+(2**8)*156+  0, (2**17)*0+(2**8)*168+ 93, (2**17)*0+(2**8)*171+107, (2**17)*0+(2**8)*238+ 32, (2**17)*0+(2**8)*281+109, (2**17)*1+(2**8)*320+ 43, 
(2**17)*0+(2**8)* 13+  0, (2**17)*0+(2**8)* 15+ 49, (2**17)*0+(2**8)* 15+121, (2**17)*0+(2**8)* 20+ 46, (2**17)*0+(2**8)* 29+165, (2**17)*0+(2**8)* 31+  0, (2**17)*0+(2**8)* 45+156, (2**17)*0+(2**8)* 49+  0, (2**17)*0+(2**8)* 57+117, (2**17)*0+(2**8)* 67+  0, (2**17)*0+(2**8)* 85+  0, (2**17)*0+(2**8)*103+  0, (2**17)*0+(2**8)*117+ 85, (2**17)*0+(2**8)*121+  0, (2**17)*0+(2**8)*136+143, (2**17)*0+(2**8)*139+  0, (2**17)*0+(2**8)*145+ 34, (2**17)*0+(2**8)*157+  0, (2**17)*0+(2**8)*162+156, (2**17)*0+(2**8)*205+101, (2**17)*0+(2**8)*231+ 31, (2**17)*0+(2**8)*244+ 44, (2**17)*0+(2**8)*247+149, (2**17)*0+(2**8)*263+ 26, (2**17)*0+(2**8)*265+ 54, (2**17)*0+(2**8)*287+122, (2**17)*0+(2**8)*300+ 18, (2**17)*1+(2**8)*319+157, 
(2**17)*0+(2**8)*  6+ 62, (2**17)*0+(2**8)* 10+115, (2**17)*0+(2**8)* 14+  0, (2**17)*0+(2**8)* 19+121, (2**17)*0+(2**8)* 32+  0, (2**17)*0+(2**8)* 50+  0, (2**17)*0+(2**8)* 68+  0, (2**17)*0+(2**8)* 75+144, (2**17)*0+(2**8)* 81+166, (2**17)*0+(2**8)* 86+  0, (2**17)*0+(2**8)*104+  0, (2**17)*0+(2**8)*113+ 33, (2**17)*0+(2**8)*122+  0, (2**17)*0+(2**8)*122+ 97, (2**17)*0+(2**8)*127+142, (2**17)*0+(2**8)*140+  0, (2**17)*0+(2**8)*158+  0, (2**17)*0+(2**8)*165+113, (2**17)*0+(2**8)*183+129, (2**17)*0+(2**8)*203+ 80, (2**17)*0+(2**8)*210+ 51, (2**17)*0+(2**8)*227+119, (2**17)*0+(2**8)*232+175, (2**17)*0+(2**8)*257+134, (2**17)*0+(2**8)*261+ 21, (2**17)*0+(2**8)*304+ 82, (2**17)*0+(2**8)*309+ 20, (2**17)*1+(2**8)*315+157, 
(2**17)*0+(2**8)* 13+168, (2**17)*0+(2**8)* 15+  0, (2**17)*0+(2**8)* 17+140, (2**17)*0+(2**8)* 33+  0, (2**17)*0+(2**8)* 51+  0, (2**17)*0+(2**8)* 66+ 10, (2**17)*0+(2**8)* 69+  0, (2**17)*0+(2**8)* 83+122, (2**17)*0+(2**8)* 85+110, (2**17)*0+(2**8)* 87+  0, (2**17)*0+(2**8)* 99+ 58, (2**17)*0+(2**8)*105+  0, (2**17)*0+(2**8)*123+  0, (2**17)*0+(2**8)*129+ 69, (2**17)*0+(2**8)*141+  0, (2**17)*0+(2**8)*151+ 73, (2**17)*0+(2**8)*159+  0, (2**17)*0+(2**8)*164+ 69, (2**17)*0+(2**8)*184+109, (2**17)*0+(2**8)*190+ 26, (2**17)*0+(2**8)*211+ 47, (2**17)*0+(2**8)*211+ 62, (2**17)*0+(2**8)*225+ 87, (2**17)*0+(2**8)*266+ 40, (2**17)*0+(2**8)*274+ 78, (2**17)*0+(2**8)*277+147, (2**17)*0+(2**8)*290+159, (2**17)*1+(2**8)*317+ 99, 
(2**17)*0+(2**8)* 16+  0, (2**17)*0+(2**8)* 33+172, (2**17)*0+(2**8)* 34+  0, (2**17)*0+(2**8)* 37+ 80, (2**17)*0+(2**8)* 52+  0, (2**17)*0+(2**8)* 59+ 88, (2**17)*0+(2**8)* 70+  0, (2**17)*0+(2**8)* 88+  0, (2**17)*0+(2**8)* 98+115, (2**17)*0+(2**8)*106+  0, (2**17)*0+(2**8)*124+  0, (2**17)*0+(2**8)*125+113, (2**17)*0+(2**8)*142+  0, (2**17)*0+(2**8)*149+ 36, (2**17)*0+(2**8)*160+  0, (2**17)*0+(2**8)*166+ 81, (2**17)*0+(2**8)*171+ 43, (2**17)*0+(2**8)*176+150, (2**17)*0+(2**8)*180+170, (2**17)*0+(2**8)*215+160, (2**17)*0+(2**8)*227+159, (2**17)*0+(2**8)*238+123, (2**17)*0+(2**8)*239+ 89, (2**17)*0+(2**8)*265+139, (2**17)*0+(2**8)*273+159, (2**17)*0+(2**8)*289+ 30, (2**17)*0+(2**8)*304+ 18, (2**17)*1+(2**8)*312+ 71, 
(2**17)*0+(2**8)*  3+118, (2**17)*0+(2**8)* 10+154, (2**17)*0+(2**8)* 13+ 39, (2**17)*0+(2**8)* 17+  0, (2**17)*0+(2**8)* 35+  0, (2**17)*0+(2**8)* 50+ 12, (2**17)*0+(2**8)* 53+  0, (2**17)*0+(2**8)* 54+ 72, (2**17)*0+(2**8)* 71+  0, (2**17)*0+(2**8)* 71+ 40, (2**17)*0+(2**8)* 89+  0, (2**17)*0+(2**8)* 89+113, (2**17)*0+(2**8)*107+  0, (2**17)*0+(2**8)*125+  0, (2**17)*0+(2**8)*133+ 36, (2**17)*0+(2**8)*141+ 16, (2**17)*0+(2**8)*143+  0, (2**17)*0+(2**8)*156+ 99, (2**17)*0+(2**8)*157+129, (2**17)*0+(2**8)*161+  0, (2**17)*0+(2**8)*187+168, (2**17)*0+(2**8)*187+ 19, (2**17)*0+(2**8)*201+155, (2**17)*0+(2**8)*248+ 53, (2**17)*0+(2**8)*256+165, (2**17)*0+(2**8)*258+ 41, (2**17)*0+(2**8)*279+ 69, (2**17)*1+(2**8)*285+ 12, 
(2**17)*0+(2**8)* 35+ 60, (2**17)*0+(2**8)* 64+145, (2**17)*0+(2**8)* 86+ 51, (2**17)*0+(2**8)* 97+118, (2**17)*0+(2**8)*153+ 32, (2**17)*0+(2**8)*162+  0, (2**17)*0+(2**8)*163+145, (2**17)*0+(2**8)*173+150, (2**17)*0+(2**8)*175+ 98, (2**17)*0+(2**8)*180+  0, (2**17)*0+(2**8)*188+156, (2**17)*0+(2**8)*198+  0, (2**17)*0+(2**8)*199+104, (2**17)*0+(2**8)*215+ 63, (2**17)*0+(2**8)*216+  0, (2**17)*0+(2**8)*219+ 57, (2**17)*0+(2**8)*234+  0, (2**17)*0+(2**8)*246+ 37, (2**17)*0+(2**8)*252+  0, (2**17)*0+(2**8)*253+  4, (2**17)*0+(2**8)*270+  0, (2**17)*0+(2**8)*274+174, (2**17)*0+(2**8)*286+108, (2**17)*0+(2**8)*288+  0, (2**17)*0+(2**8)*288+ 47, (2**17)*0+(2**8)*293+ 29, (2**17)*0+(2**8)*306+  0, (2**17)*1+(2**8)*316+ 32, 
(2**17)*0+(2**8)* 30+130, (2**17)*0+(2**8)* 44+140, (2**17)*0+(2**8)* 56+117, (2**17)*0+(2**8)* 62+ 86, (2**17)*0+(2**8)* 94+ 51, (2**17)*0+(2**8)*144+160, (2**17)*0+(2**8)*163+  0, (2**17)*0+(2**8)*165+174, (2**17)*0+(2**8)*169+ 94, (2**17)*0+(2**8)*174+148, (2**17)*0+(2**8)*181+  0, (2**17)*0+(2**8)*193+164, (2**17)*0+(2**8)*199+  0, (2**17)*0+(2**8)*206+ 40, (2**17)*0+(2**8)*217+  0, (2**17)*0+(2**8)*235+  0, (2**17)*0+(2**8)*237+ 15, (2**17)*0+(2**8)*249+100, (2**17)*0+(2**8)*253+  0, (2**17)*0+(2**8)*262+107, (2**17)*0+(2**8)*271+  0, (2**17)*0+(2**8)*280+148, (2**17)*0+(2**8)*281+ 18, (2**17)*0+(2**8)*289+  0, (2**17)*0+(2**8)*302+ 18, (2**17)*0+(2**8)*305+117, (2**17)*0+(2**8)*307+  0, (2**17)*1+(2**8)*320+150, 
(2**17)*0+(2**8)*  0+ 80, (2**17)*0+(2**8)*  8+  6, (2**17)*0+(2**8)* 27+ 58, (2**17)*0+(2**8)* 34+ 96, (2**17)*0+(2**8)* 36+ 24, (2**17)*0+(2**8)* 40+ 94, (2**17)*0+(2**8)* 62+ 26, (2**17)*0+(2**8)* 79+114, (2**17)*0+(2**8)* 82+121, (2**17)*0+(2**8)*109+144, (2**17)*0+(2**8)*164+  0, (2**17)*0+(2**8)*178+ 37, (2**17)*0+(2**8)*182+  0, (2**17)*0+(2**8)*200+  0, (2**17)*0+(2**8)*218+  0, (2**17)*0+(2**8)*220+119, (2**17)*0+(2**8)*236+  0, (2**17)*0+(2**8)*254+  0, (2**17)*0+(2**8)*260+ 56, (2**17)*0+(2**8)*262+103, (2**17)*0+(2**8)*272+  0, (2**17)*0+(2**8)*286+153, (2**17)*0+(2**8)*290+  0, (2**17)*0+(2**8)*299+130, (2**17)*0+(2**8)*305+ 40, (2**17)*0+(2**8)*308+  0, (2**17)*0+(2**8)*308+ 42, (2**17)*1+(2**8)*321+141, 
(2**17)*0+(2**8)* 12+ 33, (2**17)*0+(2**8)* 16+ 59, (2**17)*0+(2**8)* 20+ 94, (2**17)*0+(2**8)* 23+ 47, (2**17)*0+(2**8)* 52+ 18, (2**17)*0+(2**8)* 69+ 89, (2**17)*0+(2**8)* 78+ 14, (2**17)*0+(2**8)*106+129, (2**17)*0+(2**8)*110+154, (2**17)*0+(2**8)*138+ 84, (2**17)*0+(2**8)*146+ 61, (2**17)*0+(2**8)*152+ 37, (2**17)*0+(2**8)*165+  0, (2**17)*0+(2**8)*167+ 92, (2**17)*0+(2**8)*183+  0, (2**17)*0+(2**8)*201+  0, (2**17)*0+(2**8)*201+ 95, (2**17)*0+(2**8)*219+  0, (2**17)*0+(2**8)*233+ 25, (2**17)*0+(2**8)*237+  0, (2**17)*0+(2**8)*241+ 30, (2**17)*0+(2**8)*255+  0, (2**17)*0+(2**8)*267+ 35, (2**17)*0+(2**8)*270+ 88, (2**17)*0+(2**8)*273+  0, (2**17)*0+(2**8)*291+  0, (2**17)*0+(2**8)*297+101, (2**17)*1+(2**8)*309+  0, 
(2**17)*0+(2**8)*  4+156, (2**17)*0+(2**8)*  5+ 60, (2**17)*0+(2**8)* 22+ 37, (2**17)*0+(2**8)* 24+ 79, (2**17)*0+(2**8)* 45+ 16, (2**17)*0+(2**8)* 61+ 32, (2**17)*0+(2**8)* 77+ 80, (2**17)*0+(2**8)* 80+ 64, (2**17)*0+(2**8)*115+111, (2**17)*0+(2**8)*152+138, (2**17)*0+(2**8)*166+  0, (2**17)*0+(2**8)*176+ 41, (2**17)*0+(2**8)*184+  0, (2**17)*0+(2**8)*202+  0, (2**17)*0+(2**8)*213+ 64, (2**17)*0+(2**8)*220+  0, (2**17)*0+(2**8)*230+123, (2**17)*0+(2**8)*238+  0, (2**17)*0+(2**8)*252+ 49, (2**17)*0+(2**8)*252+ 90, (2**17)*0+(2**8)*256+  0, (2**17)*0+(2**8)*274+  0, (2**17)*0+(2**8)*276+ 90, (2**17)*0+(2**8)*288+162, (2**17)*0+(2**8)*292+  0, (2**17)*0+(2**8)*296+ 97, (2**17)*0+(2**8)*310+  0, (2**17)*1+(2**8)*317+149, 
(2**17)*0+(2**8)*  8+ 72, (2**17)*0+(2**8)* 16+115, (2**17)*0+(2**8)* 59+153, (2**17)*0+(2**8)* 61+  3, (2**17)*0+(2**8)*121+105, (2**17)*0+(2**8)*122+ 86, (2**17)*0+(2**8)*132+175, (2**17)*0+(2**8)*133+155, (2**17)*0+(2**8)*159+ 74, (2**17)*0+(2**8)*167+  0, (2**17)*0+(2**8)*173+ 82, (2**17)*0+(2**8)*180+150, (2**17)*0+(2**8)*185+  0, (2**17)*0+(2**8)*194+119, (2**17)*0+(2**8)*203+  0, (2**17)*0+(2**8)*208+150, (2**17)*0+(2**8)*208+ 13, (2**17)*0+(2**8)*221+  0, (2**17)*0+(2**8)*236+123, (2**17)*0+(2**8)*236+121, (2**17)*0+(2**8)*239+  0, (2**17)*0+(2**8)*254+ 44, (2**17)*0+(2**8)*257+  0, (2**17)*0+(2**8)*267+  8, (2**17)*0+(2**8)*275+  0, (2**17)*0+(2**8)*293+  0, (2**17)*0+(2**8)*311+  0, (2**17)*1+(2**8)*311+ 42, 
(2**17)*0+(2**8)* 40+ 98, (2**17)*0+(2**8)* 60+126, (2**17)*0+(2**8)* 78+ 75, (2**17)*0+(2**8)* 87+159, (2**17)*0+(2**8)*113+ 72, (2**17)*0+(2**8)*121+139, (2**17)*0+(2**8)*135+ 97, (2**17)*0+(2**8)*139+ 72, (2**17)*0+(2**8)*151+146, (2**17)*0+(2**8)*164+ 23, (2**17)*0+(2**8)*167+ 48, (2**17)*0+(2**8)*168+  0, (2**17)*0+(2**8)*170+148, (2**17)*0+(2**8)*181+ 83, (2**17)*0+(2**8)*183+154, (2**17)*0+(2**8)*186+  0, (2**17)*0+(2**8)*204+  0, (2**17)*0+(2**8)*214+ 31, (2**17)*0+(2**8)*222+  0, (2**17)*0+(2**8)*230+ 25, (2**17)*0+(2**8)*240+  0, (2**17)*0+(2**8)*255+143, (2**17)*0+(2**8)*257+ 75, (2**17)*0+(2**8)*258+  0, (2**17)*0+(2**8)*276+  0, (2**17)*0+(2**8)*294+  0, (2**17)*0+(2**8)*310+107, (2**17)*1+(2**8)*312+  0, 
(2**17)*0+(2**8)*  1+133, (2**17)*0+(2**8)*  7+ 60, (2**17)*0+(2**8)* 24+150, (2**17)*0+(2**8)* 28+136, (2**17)*0+(2**8)* 36+115, (2**17)*0+(2**8)* 58+ 97, (2**17)*0+(2**8)* 81+155, (2**17)*0+(2**8)* 91+ 59, (2**17)*0+(2**8)*116+ 62, (2**17)*0+(2**8)*136+ 63, (2**17)*0+(2**8)*162+ 71, (2**17)*0+(2**8)*169+  0, (2**17)*0+(2**8)*187+  0, (2**17)*0+(2**8)*203+153, (2**17)*0+(2**8)*205+  0, (2**17)*0+(2**8)*218+ 34, (2**17)*0+(2**8)*223+  0, (2**17)*0+(2**8)*241+  0, (2**17)*0+(2**8)*246+171, (2**17)*0+(2**8)*254+119, (2**17)*0+(2**8)*259+  0, (2**17)*0+(2**8)*277+  0, (2**17)*0+(2**8)*278+ 85, (2**17)*0+(2**8)*295+  0, (2**17)*0+(2**8)*296+ 36, (2**17)*0+(2**8)*310+143, (2**17)*0+(2**8)*313+  0, (2**17)*1+(2**8)*318+ 39, 
(2**17)*0+(2**8)*  6+157, (2**17)*0+(2**8)* 11+121, (2**17)*0+(2**8)* 26+ 71, (2**17)*0+(2**8)* 30+ 39, (2**17)*0+(2**8)* 47+144, (2**17)*0+(2**8)* 55+ 21, (2**17)*0+(2**8)* 88+ 90, (2**17)*0+(2**8)*102+170, (2**17)*0+(2**8)*109+ 58, (2**17)*0+(2**8)*150+ 87, (2**17)*0+(2**8)*170+  0, (2**17)*0+(2**8)*179+  7, (2**17)*0+(2**8)*188+  0, (2**17)*0+(2**8)*206+  0, (2**17)*0+(2**8)*209+131, (2**17)*0+(2**8)*224+  0, (2**17)*0+(2**8)*225+ 30, (2**17)*0+(2**8)*242+  0, (2**17)*0+(2**8)*250+168, (2**17)*0+(2**8)*260+  0, (2**17)*0+(2**8)*269+177, (2**17)*0+(2**8)*278+  0, (2**17)*0+(2**8)*280+ 33, (2**17)*0+(2**8)*293+ 41, (2**17)*0+(2**8)*296+  0, (2**17)*0+(2**8)*303+173, (2**17)*0+(2**8)*314+  0, (2**17)*1+(2**8)*323+ 94, 
(2**17)*0+(2**8)*  9+ 48, (2**17)*0+(2**8)* 15+106, (2**17)*0+(2**8)* 27+ 32, (2**17)*0+(2**8)* 42+ 47, (2**17)*0+(2**8)* 60+ 53, (2**17)*0+(2**8)* 70+ 71, (2**17)*0+(2**8)* 72+ 23, (2**17)*0+(2**8)* 80+166, (2**17)*0+(2**8)*123+132, (2**17)*0+(2**8)*140+ 90, (2**17)*0+(2**8)*145+ 66, (2**17)*0+(2**8)*160+ 48, (2**17)*0+(2**8)*164+  2, (2**17)*0+(2**8)*171+  0, (2**17)*0+(2**8)*185+  3, (2**17)*0+(2**8)*189+  0, (2**17)*0+(2**8)*205+ 21, (2**17)*0+(2**8)*207+  0, (2**17)*0+(2**8)*225+  0, (2**17)*0+(2**8)*243+  0, (2**17)*0+(2**8)*259+ 19, (2**17)*0+(2**8)*261+  0, (2**17)*0+(2**8)*268+165, (2**17)*0+(2**8)*279+  0, (2**17)*0+(2**8)*282+127, (2**17)*0+(2**8)*290+171, (2**17)*0+(2**8)*297+  0, (2**17)*1+(2**8)*315+  0, 
(2**17)*0+(2**8)* 14+ 29, (2**17)*0+(2**8)* 17+ 65, (2**17)*0+(2**8)* 51+ 85, (2**17)*0+(2**8)* 93+ 34, (2**17)*0+(2**8)*104+142, (2**17)*0+(2**8)*160+  8, (2**17)*0+(2**8)*172+  0, (2**17)*0+(2**8)*172+ 87, (2**17)*0+(2**8)*190+  0, (2**17)*0+(2**8)*194+ 51, (2**17)*0+(2**8)*195+149, (2**17)*0+(2**8)*200+ 24, (2**17)*0+(2**8)*208+  0, (2**17)*0+(2**8)*216+163, (2**17)*0+(2**8)*226+  0, (2**17)*0+(2**8)*229+ 77, (2**17)*0+(2**8)*235+110, (2**17)*0+(2**8)*244+  0, (2**17)*0+(2**8)*251+ 92, (2**17)*0+(2**8)*262+  0, (2**17)*0+(2**8)*270+130, (2**17)*0+(2**8)*276+ 28, (2**17)*0+(2**8)*280+  0, (2**17)*0+(2**8)*294+112, (2**17)*0+(2**8)*298+  0, (2**17)*0+(2**8)*301+ 78, (2**17)*0+(2**8)*316+  0, (2**17)*1+(2**8)*316+121, 
(2**17)*0+(2**8)* 29+ 62, (2**17)*0+(2**8)* 38+ 77, (2**17)*0+(2**8)* 73+113, (2**17)*0+(2**8)*111+ 48, (2**17)*0+(2**8)*130+ 61, (2**17)*0+(2**8)*137+106, (2**17)*0+(2**8)*147+155, (2**17)*0+(2**8)*163+ 87, (2**17)*0+(2**8)*166+ 29, (2**17)*0+(2**8)*173+  0, (2**17)*0+(2**8)*174+ 88, (2**17)*0+(2**8)*191+  0, (2**17)*0+(2**8)*196+ 49, (2**17)*0+(2**8)*209+  0, (2**17)*0+(2**8)*210+  4, (2**17)*0+(2**8)*217+ 93, (2**17)*0+(2**8)*227+  0, (2**17)*0+(2**8)*229+  5, (2**17)*0+(2**8)*234+124, (2**17)*0+(2**8)*245+  0, (2**17)*0+(2**8)*263+  0, (2**17)*0+(2**8)*263+142, (2**17)*0+(2**8)*264+ 92, (2**17)*0+(2**8)*281+  0, (2**17)*0+(2**8)*282+105, (2**17)*0+(2**8)*299+  0, (2**17)*0+(2**8)*317+  0, (2**17)*1+(2**8)*323+ 55, 
(2**17)*0+(2**8)*  6+ 92, (2**17)*0+(2**8)*  9+106, (2**17)*0+(2**8)* 76+ 31, (2**17)*0+(2**8)*119+108, (2**17)*0+(2**8)*158+ 42, (2**17)*0+(2**8)*169+ 15, (2**17)*0+(2**8)*174+  0, (2**17)*0+(2**8)*192+  0, (2**17)*0+(2**8)*193+ 13, (2**17)*0+(2**8)*197+ 89, (2**17)*0+(2**8)*204+ 14, (2**17)*0+(2**8)*210+  0, (2**17)*0+(2**8)*212+ 32, (2**17)*0+(2**8)*226+123, (2**17)*0+(2**8)*228+  0, (2**17)*0+(2**8)*228+ 98, (2**17)*0+(2**8)*245+ 27, (2**17)*0+(2**8)*246+  0, (2**17)*0+(2**8)*258+ 93, (2**17)*0+(2**8)*264+  0, (2**17)*0+(2**8)*269+126, (2**17)*0+(2**8)*272+177, (2**17)*0+(2**8)*282+  0, (2**17)*0+(2**8)*291+ 98, (2**17)*0+(2**8)*292+176, (2**17)*0+(2**8)*300+  0, (2**17)*0+(2**8)*306+ 44, (2**17)*1+(2**8)*318+  0, 
(2**17)*0+(2**8)*  0+155, (2**17)*0+(2**8)* 43+100, (2**17)*0+(2**8)* 69+ 30, (2**17)*0+(2**8)* 82+ 43, (2**17)*0+(2**8)* 85+148, (2**17)*0+(2**8)*101+ 25, (2**17)*0+(2**8)*103+ 53, (2**17)*0+(2**8)*125+121, (2**17)*0+(2**8)*138+ 17, (2**17)*0+(2**8)*157+156, (2**17)*0+(2**8)*175+  0, (2**17)*0+(2**8)*177+ 49, (2**17)*0+(2**8)*177+121, (2**17)*0+(2**8)*182+ 46, (2**17)*0+(2**8)*191+165, (2**17)*0+(2**8)*193+  0, (2**17)*0+(2**8)*207+156, (2**17)*0+(2**8)*211+  0, (2**17)*0+(2**8)*219+117, (2**17)*0+(2**8)*229+  0, (2**17)*0+(2**8)*247+  0, (2**17)*0+(2**8)*265+  0, (2**17)*0+(2**8)*279+ 85, (2**17)*0+(2**8)*283+  0, (2**17)*0+(2**8)*298+143, (2**17)*0+(2**8)*301+  0, (2**17)*0+(2**8)*307+ 34, (2**17)*1+(2**8)*319+  0, 
(2**17)*0+(2**8)*  3+112, (2**17)*0+(2**8)* 21+128, (2**17)*0+(2**8)* 41+ 79, (2**17)*0+(2**8)* 48+ 50, (2**17)*0+(2**8)* 65+118, (2**17)*0+(2**8)* 70+174, (2**17)*0+(2**8)* 95+133, (2**17)*0+(2**8)* 99+ 20, (2**17)*0+(2**8)*142+ 81, (2**17)*0+(2**8)*147+ 19, (2**17)*0+(2**8)*153+156, (2**17)*0+(2**8)*168+ 62, (2**17)*0+(2**8)*172+115, (2**17)*0+(2**8)*176+  0, (2**17)*0+(2**8)*181+121, (2**17)*0+(2**8)*194+  0, (2**17)*0+(2**8)*212+  0, (2**17)*0+(2**8)*230+  0, (2**17)*0+(2**8)*237+144, (2**17)*0+(2**8)*243+166, (2**17)*0+(2**8)*248+  0, (2**17)*0+(2**8)*266+  0, (2**17)*0+(2**8)*275+ 33, (2**17)*0+(2**8)*284+  0, (2**17)*0+(2**8)*284+ 97, (2**17)*0+(2**8)*289+142, (2**17)*0+(2**8)*302+  0, (2**17)*1+(2**8)*320+  0, 
(2**17)*0+(2**8)*  2+ 68, (2**17)*0+(2**8)* 22+108, (2**17)*0+(2**8)* 28+ 25, (2**17)*0+(2**8)* 49+ 46, (2**17)*0+(2**8)* 49+ 61, (2**17)*0+(2**8)* 63+ 86, (2**17)*0+(2**8)*104+ 39, (2**17)*0+(2**8)*112+ 77, (2**17)*0+(2**8)*115+146, (2**17)*0+(2**8)*128+158, (2**17)*0+(2**8)*155+ 98, (2**17)*0+(2**8)*175+168, (2**17)*0+(2**8)*177+  0, (2**17)*0+(2**8)*179+140, (2**17)*0+(2**8)*195+  0, (2**17)*0+(2**8)*213+  0, (2**17)*0+(2**8)*228+ 10, (2**17)*0+(2**8)*231+  0, (2**17)*0+(2**8)*245+122, (2**17)*0+(2**8)*247+110, (2**17)*0+(2**8)*249+  0, (2**17)*0+(2**8)*261+ 58, (2**17)*0+(2**8)*267+  0, (2**17)*0+(2**8)*285+  0, (2**17)*0+(2**8)*291+ 69, (2**17)*0+(2**8)*303+  0, (2**17)*0+(2**8)*313+ 73, (2**17)*1+(2**8)*321+  0, 
(2**17)*0+(2**8)*  4+ 80, (2**17)*0+(2**8)*  9+ 42, (2**17)*0+(2**8)* 14+149, (2**17)*0+(2**8)* 18+169, (2**17)*0+(2**8)* 53+159, (2**17)*0+(2**8)* 65+158, (2**17)*0+(2**8)* 76+122, (2**17)*0+(2**8)* 77+ 88, (2**17)*0+(2**8)*103+138, (2**17)*0+(2**8)*111+158, (2**17)*0+(2**8)*127+ 29, (2**17)*0+(2**8)*142+ 17, (2**17)*0+(2**8)*150+ 70, (2**17)*0+(2**8)*178+  0, (2**17)*0+(2**8)*195+172, (2**17)*0+(2**8)*196+  0, (2**17)*0+(2**8)*199+ 80, (2**17)*0+(2**8)*214+  0, (2**17)*0+(2**8)*221+ 88, (2**17)*0+(2**8)*232+  0, (2**17)*0+(2**8)*250+  0, (2**17)*0+(2**8)*260+115, (2**17)*0+(2**8)*268+  0, (2**17)*0+(2**8)*286+  0, (2**17)*0+(2**8)*287+113, (2**17)*0+(2**8)*304+  0, (2**17)*0+(2**8)*311+ 36, (2**17)*1+(2**8)*322+  0, 
(2**17)*0+(2**8)* 25+167, (2**17)*0+(2**8)* 25+ 18, (2**17)*0+(2**8)* 39+154, (2**17)*0+(2**8)* 86+ 52, (2**17)*0+(2**8)* 94+164, (2**17)*0+(2**8)* 96+ 40, (2**17)*0+(2**8)*117+ 68, (2**17)*0+(2**8)*123+ 11, (2**17)*0+(2**8)*165+118, (2**17)*0+(2**8)*172+154, (2**17)*0+(2**8)*175+ 39, (2**17)*0+(2**8)*179+  0, (2**17)*0+(2**8)*197+  0, (2**17)*0+(2**8)*212+ 12, (2**17)*0+(2**8)*215+  0, (2**17)*0+(2**8)*216+ 72, (2**17)*0+(2**8)*233+  0, (2**17)*0+(2**8)*233+ 40, (2**17)*0+(2**8)*251+  0, (2**17)*0+(2**8)*251+113, (2**17)*0+(2**8)*269+  0, (2**17)*0+(2**8)*287+  0, (2**17)*0+(2**8)*295+ 36, (2**17)*0+(2**8)*303+ 16, (2**17)*0+(2**8)*305+  0, (2**17)*0+(2**8)*318+ 99, (2**17)*0+(2**8)*319+129, (2**17)*1+(2**8)*323+  0);


begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector(EdgeMapMemory(conv_integer(Addr)),18);
		end if;
	end process;
end Behavioral;
