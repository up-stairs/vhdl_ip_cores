LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CNP_Output_Edge_Memory is
	Port (
		clk			: in  std_logic;

		RdAddr		: in  std_logic_vector(13 downto 0);
		Do			: out std_logic_vector(16 downto 0)
	);
end CNP_Output_Edge_Memory;

architecture Behavioral of CNP_Output_Edge_Memory is
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 11672-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
  14*2048+  24,   45*2048+  25,   45*2048+  26, 
  32*2048+  51,   45*2048+  52,   45*2048+  53, 
  11*2048+  54,   45*2048+  55,   45*2048+  56, 
  28*2048+  57,   45*2048+  58,   45*2048+  59, 
  27*2048+  76,   45*2048+  77,   45*2048+  78, 
  32*2048+  99,   45*2048+ 100,   45*2048+ 101, 
  18*2048+ 102,   45*2048+ 103,   45*2048+ 104, 
  40*2048+ 105,   45*2048+ 106,   45*2048+ 107, 
   8*2048+ 112,   45*2048+ 113,   45*2048+ 114, 
  14*2048+ 159,   45*2048+ 160,   45*2048+ 161, 
  32*2048+ 186,   45*2048+ 187,   45*2048+ 188, 
  11*2048+ 189,   45*2048+ 190,   45*2048+ 191, 
  28*2048+ 192,   45*2048+ 193,   45*2048+ 194, 
  27*2048+ 211,   45*2048+ 212,   45*2048+ 213, 
  32*2048+ 234,   45*2048+ 235,   45*2048+ 236, 
  18*2048+ 237,   45*2048+ 238,   45*2048+ 239, 
  40*2048+ 240,   45*2048+ 241,   45*2048+ 242, 
   8*2048+ 247,   45*2048+ 248,   45*2048+ 249, 
  15*2048+ 294,   45*2048+ 295,   45*2048+ 296, 
  32*2048+ 321,   45*2048+ 322,   45*2048+ 323, 
  11*2048+ 324,   45*2048+ 325,   45*2048+ 326, 
  28*2048+ 327,   45*2048+ 328,   45*2048+ 329, 
  28*2048+ 346,   45*2048+ 347,   45*2048+ 348, 
  32*2048+ 369,   45*2048+ 370,   45*2048+ 371, 
  18*2048+ 372,   45*2048+ 373,   45*2048+ 374, 
  40*2048+ 375,   45*2048+ 376,   45*2048+ 377, 
   8*2048+ 382,   45*2048+ 383,   45*2048+ 384, 
  15*2048+ 429,   45*2048+ 430,   45*2048+ 431, 
  32*2048+ 456,   45*2048+ 457,   45*2048+ 458, 
  12*2048+ 459,   45*2048+ 460,   45*2048+ 461, 
  28*2048+ 462,   45*2048+ 463,   45*2048+ 464, 
  28*2048+ 481,   45*2048+ 482,   45*2048+ 483, 
  32*2048+ 504,   45*2048+ 505,   45*2048+ 506, 
  18*2048+ 507,   45*2048+ 508,   45*2048+ 509, 
  40*2048+ 510,   45*2048+ 511,   45*2048+ 512, 
   8*2048+ 517,   45*2048+ 518,   45*2048+ 519, 
  15*2048+ 564,   45*2048+ 565,   45*2048+ 566, 
  33*2048+ 591,   45*2048+ 592,   45*2048+ 593, 
  12*2048+ 594,   45*2048+ 595,   45*2048+ 596, 
  28*2048+ 597,   45*2048+ 598,   45*2048+ 599, 
  28*2048+ 616,   45*2048+ 617,   45*2048+ 618, 
  32*2048+ 639,   45*2048+ 640,   45*2048+ 641, 
  18*2048+ 642,   45*2048+ 643,   45*2048+ 644, 
  40*2048+ 645,   45*2048+ 646,   45*2048+ 647, 
   8*2048+ 652,   45*2048+ 653,   45*2048+ 654, 
  15*2048+ 699,   45*2048+ 700,   45*2048+ 701, 
  33*2048+ 726,   45*2048+ 727,   45*2048+ 728, 
  12*2048+ 729,   45*2048+ 730,   45*2048+ 731, 
  28*2048+ 732,   45*2048+ 733,   45*2048+ 734, 
  28*2048+ 751,   45*2048+ 752,   45*2048+ 753, 
  32*2048+ 774,   45*2048+ 775,   45*2048+ 776, 
  19*2048+ 777,   45*2048+ 778,   45*2048+ 779, 
  41*2048+ 780,   45*2048+ 781,   45*2048+ 782, 
   8*2048+ 787,   45*2048+ 788,   45*2048+ 789, 
  15*2048+ 834,   45*2048+ 835,   45*2048+ 836, 
  33*2048+ 861,   45*2048+ 862,   45*2048+ 863, 
  12*2048+ 864,   45*2048+ 865,   45*2048+ 866, 
  29*2048+ 867,   45*2048+ 868,   45*2048+ 869, 
  28*2048+ 886,   45*2048+ 887,   45*2048+ 888, 
  32*2048+ 909,   45*2048+ 910,   45*2048+ 911, 
  19*2048+ 912,   45*2048+ 913,   45*2048+ 914, 
  41*2048+ 915,   45*2048+ 916,   45*2048+ 917, 
   8*2048+ 922,   45*2048+ 923,   45*2048+ 924, 
  15*2048+ 969,   45*2048+ 970,   45*2048+ 971, 
  33*2048+ 996,   45*2048+ 997,   45*2048+ 998, 
  12*2048+ 999,   45*2048+1000,   45*2048+1001, 
  29*2048+1002,   45*2048+1003,   45*2048+1004, 
  28*2048+1021,   45*2048+1022,   45*2048+1023, 
  33*2048+1044,   45*2048+1045,   45*2048+1046, 
  19*2048+1047,   45*2048+1048,   45*2048+1049, 
  41*2048+1050,   45*2048+1051,   45*2048+1052, 
   9*2048+1057,   45*2048+1058,   45*2048+1059, 
  32*2048+   0,   44*2048+   1,   45*2048+   2,   44*2048+   3, 
  33*2048+   4,   21*2048+   5,   45*2048+   6,   45*2048+   7, 
   6*2048+   8,   32*2048+   9,   45*2048+  10,   45*2048+  11, 
  19*2048+  12,   36*2048+  13,   45*2048+  14,   45*2048+  15, 
  39*2048+  16,   27*2048+  17,   45*2048+  18,   45*2048+  19, 
  17*2048+  20,   24*2048+  21,   45*2048+  22,   45*2048+  23, 
   6*2048+  27,   31*2048+  28,   45*2048+  29,   45*2048+  30, 
  30*2048+  31,   18*2048+  32,   45*2048+  33,   45*2048+  34, 
   7*2048+  35,   27*2048+  36,   45*2048+  37,   45*2048+  38, 
   7*2048+  39,   35*2048+  40,   45*2048+  41,   45*2048+  42, 
  23*2048+  43,   34*2048+  44,   45*2048+  45,   45*2048+  46, 
  28*2048+  47,   10*2048+  48,   45*2048+  49,   45*2048+  50, 
  44*2048+  60,   16*2048+  61,   45*2048+  62,   45*2048+  63, 
   9*2048+  64,    6*2048+  65,   45*2048+  66,   45*2048+  67, 
   7*2048+  68,    0*2048+  69,   45*2048+  70,   45*2048+  71, 
  18*2048+  72,   34*2048+  73,   45*2048+  74,   45*2048+  75, 
  32*2048+  79,    8*2048+  80,   45*2048+  81,   45*2048+  82, 
   3*2048+  83,   33*2048+  84,   45*2048+  85,   45*2048+  86, 
  25*2048+  87,   25*2048+  88,   45*2048+  89,   45*2048+  90, 
  27*2048+  91,   24*2048+  92,   45*2048+  93,   45*2048+  94, 
   2*2048+  95,    3*2048+  96,   45*2048+  97,   45*2048+  98, 
  30*2048+ 108,    1*2048+ 109,   45*2048+ 110,   45*2048+ 111, 
  23*2048+ 115,   22*2048+ 116,   45*2048+ 117,   45*2048+ 118, 
   6*2048+ 119,   17*2048+ 120,   45*2048+ 121,   45*2048+ 122, 
  23*2048+ 123,   12*2048+ 124,   45*2048+ 125,   45*2048+ 126, 
  14*2048+ 127,    2*2048+ 128,   45*2048+ 129,   45*2048+ 130, 
   8*2048+ 131,   36*2048+ 132,   45*2048+ 133,   45*2048+ 134, 
  32*2048+ 135,   44*2048+ 136,   45*2048+ 137,   45*2048+ 138, 
  33*2048+ 139,   21*2048+ 140,   45*2048+ 141,   45*2048+ 142, 
  33*2048+ 143,    6*2048+ 144,   45*2048+ 145,   45*2048+ 146, 
  20*2048+ 147,   37*2048+ 148,   45*2048+ 149,   45*2048+ 150, 
  28*2048+ 151,   39*2048+ 152,   45*2048+ 153,   45*2048+ 154, 
  17*2048+ 155,   24*2048+ 156,   45*2048+ 157,   45*2048+ 158, 
   6*2048+ 162,   31*2048+ 163,   45*2048+ 164,   45*2048+ 165, 
  30*2048+ 166,   18*2048+ 167,   45*2048+ 168,   45*2048+ 169, 
   7*2048+ 170,   27*2048+ 171,   45*2048+ 172,   45*2048+ 173, 
   7*2048+ 174,   35*2048+ 175,   45*2048+ 176,   45*2048+ 177, 
  23*2048+ 178,   34*2048+ 179,   45*2048+ 180,   45*2048+ 181, 
  11*2048+ 182,   28*2048+ 183,   45*2048+ 184,   45*2048+ 185, 
  44*2048+ 195,   16*2048+ 196,   45*2048+ 197,   45*2048+ 198, 
   9*2048+ 199,    6*2048+ 200,   45*2048+ 201,   45*2048+ 202, 
   1*2048+ 203,    7*2048+ 204,   45*2048+ 205,   45*2048+ 206, 
  18*2048+ 207,   34*2048+ 208,   45*2048+ 209,   45*2048+ 210, 
  32*2048+ 214,    8*2048+ 215,   45*2048+ 216,   45*2048+ 217, 
   3*2048+ 218,   33*2048+ 219,   45*2048+ 220,   45*2048+ 221, 
  25*2048+ 222,   25*2048+ 223,   45*2048+ 224,   45*2048+ 225, 
  27*2048+ 226,   24*2048+ 227,   45*2048+ 228,   45*2048+ 229, 
   4*2048+ 230,    2*2048+ 231,   45*2048+ 232,   45*2048+ 233, 
  30*2048+ 243,    1*2048+ 244,   45*2048+ 245,   45*2048+ 246, 
  23*2048+ 250,   22*2048+ 251,   45*2048+ 252,   45*2048+ 253, 
  18*2048+ 254,    6*2048+ 255,   45*2048+ 256,   45*2048+ 257, 
  13*2048+ 258,   23*2048+ 259,   45*2048+ 260,   45*2048+ 261, 
  14*2048+ 262,    2*2048+ 263,   45*2048+ 264,   45*2048+ 265, 
   8*2048+ 266,   36*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
  32*2048+ 270,   44*2048+ 271,   45*2048+ 272,   45*2048+ 273, 
  33*2048+ 274,   21*2048+ 275,   45*2048+ 276,   45*2048+ 277, 
  33*2048+ 278,    6*2048+ 279,   45*2048+ 280,   45*2048+ 281, 
  20*2048+ 282,   37*2048+ 283,   45*2048+ 284,   45*2048+ 285, 
  28*2048+ 286,   39*2048+ 287,   45*2048+ 288,   45*2048+ 289, 
  17*2048+ 290,   24*2048+ 291,   45*2048+ 292,   45*2048+ 293, 
   6*2048+ 297,   31*2048+ 298,   45*2048+ 299,   45*2048+ 300, 
  30*2048+ 301,   18*2048+ 302,   45*2048+ 303,   45*2048+ 304, 
  28*2048+ 305,    7*2048+ 306,   45*2048+ 307,   45*2048+ 308, 
  36*2048+ 309,    7*2048+ 310,   45*2048+ 311,   45*2048+ 312, 
  23*2048+ 313,   34*2048+ 314,   45*2048+ 315,   45*2048+ 316, 
  11*2048+ 317,   28*2048+ 318,   45*2048+ 319,   45*2048+ 320, 
  44*2048+ 330,   16*2048+ 331,   45*2048+ 332,   45*2048+ 333, 
   9*2048+ 334,    6*2048+ 335,   45*2048+ 336,   45*2048+ 337, 
   1*2048+ 338,    7*2048+ 339,   45*2048+ 340,   45*2048+ 341, 
  18*2048+ 342,   34*2048+ 343,   45*2048+ 344,   45*2048+ 345, 
  33*2048+ 349,    9*2048+ 350,   45*2048+ 351,   45*2048+ 352, 
   3*2048+ 353,   33*2048+ 354,   45*2048+ 355,   45*2048+ 356, 
  26*2048+ 357,   25*2048+ 358,   45*2048+ 359,   45*2048+ 360, 
  27*2048+ 361,   24*2048+ 362,   45*2048+ 363,   45*2048+ 364, 
   4*2048+ 365,    2*2048+ 366,   45*2048+ 367,   45*2048+ 368, 
  30*2048+ 378,    1*2048+ 379,   45*2048+ 380,   45*2048+ 381, 
  23*2048+ 385,   22*2048+ 386,   45*2048+ 387,   45*2048+ 388, 
  18*2048+ 389,    6*2048+ 390,   45*2048+ 391,   45*2048+ 392, 
  13*2048+ 393,   23*2048+ 394,   45*2048+ 395,   45*2048+ 396, 
  15*2048+ 397,    3*2048+ 398,   45*2048+ 399,   45*2048+ 400, 
   8*2048+ 401,   36*2048+ 402,   45*2048+ 403,   45*2048+ 404, 
  32*2048+ 405,   44*2048+ 406,   45*2048+ 407,   45*2048+ 408, 
  33*2048+ 409,   21*2048+ 410,   45*2048+ 411,   45*2048+ 412, 
  33*2048+ 413,    6*2048+ 414,   45*2048+ 415,   45*2048+ 416, 
  20*2048+ 417,   37*2048+ 418,   45*2048+ 419,   45*2048+ 420, 
  28*2048+ 421,   39*2048+ 422,   45*2048+ 423,   45*2048+ 424, 
  17*2048+ 425,   24*2048+ 426,   45*2048+ 427,   45*2048+ 428, 
  32*2048+ 432,    6*2048+ 433,   45*2048+ 434,   45*2048+ 435, 
  30*2048+ 436,   18*2048+ 437,   45*2048+ 438,   45*2048+ 439, 
   8*2048+ 440,   28*2048+ 441,   45*2048+ 442,   45*2048+ 443, 
   8*2048+ 444,   36*2048+ 445,   45*2048+ 446,   45*2048+ 447, 
  23*2048+ 448,   34*2048+ 449,   45*2048+ 450,   45*2048+ 451, 
  11*2048+ 452,   28*2048+ 453,   45*2048+ 454,   45*2048+ 455, 
  44*2048+ 465,   16*2048+ 466,   45*2048+ 467,   45*2048+ 468, 
   9*2048+ 469,    6*2048+ 470,   45*2048+ 471,   45*2048+ 472, 
   1*2048+ 473,    7*2048+ 474,   45*2048+ 475,   45*2048+ 476, 
  18*2048+ 477,   34*2048+ 478,   45*2048+ 479,   45*2048+ 480, 
  33*2048+ 484,    9*2048+ 485,   45*2048+ 486,   45*2048+ 487, 
   3*2048+ 488,   33*2048+ 489,   45*2048+ 490,   45*2048+ 491, 
  26*2048+ 492,   25*2048+ 493,   45*2048+ 494,   45*2048+ 495, 
  27*2048+ 496,   24*2048+ 497,   45*2048+ 498,   45*2048+ 499, 
   4*2048+ 500,    2*2048+ 501,   45*2048+ 502,   45*2048+ 503, 
  30*2048+ 513,    1*2048+ 514,   45*2048+ 515,   45*2048+ 516, 
  23*2048+ 520,   22*2048+ 521,   45*2048+ 522,   45*2048+ 523, 
  18*2048+ 524,    6*2048+ 525,   45*2048+ 526,   45*2048+ 527, 
  24*2048+ 528,   13*2048+ 529,   45*2048+ 530,   45*2048+ 531, 
  15*2048+ 532,    3*2048+ 533,   45*2048+ 534,   45*2048+ 535, 
   8*2048+ 536,   36*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
  45*2048+ 540,   32*2048+ 541,   45*2048+ 542,   45*2048+ 543, 
  33*2048+ 544,   21*2048+ 545,   45*2048+ 546,   45*2048+ 547, 
   7*2048+ 548,   33*2048+ 549,   45*2048+ 550,   45*2048+ 551, 
  20*2048+ 552,   37*2048+ 553,   45*2048+ 554,   45*2048+ 555, 
  28*2048+ 556,   39*2048+ 557,   45*2048+ 558,   45*2048+ 559, 
  17*2048+ 560,   24*2048+ 561,   45*2048+ 562,   45*2048+ 563, 
  32*2048+ 567,    6*2048+ 568,   45*2048+ 569,   45*2048+ 570, 
  30*2048+ 571,   18*2048+ 572,   45*2048+ 573,   45*2048+ 574, 
   8*2048+ 575,   28*2048+ 576,   45*2048+ 577,   45*2048+ 578, 
   8*2048+ 579,   36*2048+ 580,   45*2048+ 581,   45*2048+ 582, 
  23*2048+ 583,   34*2048+ 584,   45*2048+ 585,   45*2048+ 586, 
  11*2048+ 587,   28*2048+ 588,   45*2048+ 589,   45*2048+ 590, 
  44*2048+ 600,   16*2048+ 601,   45*2048+ 602,   45*2048+ 603, 
   9*2048+ 604,    6*2048+ 605,   45*2048+ 606,   45*2048+ 607, 
   1*2048+ 608,    7*2048+ 609,   45*2048+ 610,   45*2048+ 611, 
  18*2048+ 612,   34*2048+ 613,   45*2048+ 614,   45*2048+ 615, 
  33*2048+ 619,    9*2048+ 620,   45*2048+ 621,   45*2048+ 622, 
  34*2048+ 623,    3*2048+ 624,   45*2048+ 625,   45*2048+ 626, 
  26*2048+ 627,   25*2048+ 628,   45*2048+ 629,   45*2048+ 630, 
  27*2048+ 631,   24*2048+ 632,   45*2048+ 633,   45*2048+ 634, 
   3*2048+ 635,    4*2048+ 636,   45*2048+ 637,   45*2048+ 638, 
   2*2048+ 648,   30*2048+ 649,   45*2048+ 650,   45*2048+ 651, 
  23*2048+ 655,   22*2048+ 656,   45*2048+ 657,   45*2048+ 658, 
   7*2048+ 659,   18*2048+ 660,   45*2048+ 661,   45*2048+ 662, 
  24*2048+ 663,   13*2048+ 664,   45*2048+ 665,   45*2048+ 666, 
  15*2048+ 667,    3*2048+ 668,   45*2048+ 669,   45*2048+ 670, 
   8*2048+ 671,   36*2048+ 672,   45*2048+ 673,   45*2048+ 674, 
  45*2048+ 675,   32*2048+ 676,   45*2048+ 677,   45*2048+ 678, 
  22*2048+ 679,   33*2048+ 680,   45*2048+ 681,   45*2048+ 682, 
   7*2048+ 683,   33*2048+ 684,   45*2048+ 685,   45*2048+ 686, 
  20*2048+ 687,   37*2048+ 688,   45*2048+ 689,   45*2048+ 690, 
  28*2048+ 691,   39*2048+ 692,   45*2048+ 693,   45*2048+ 694, 
  17*2048+ 695,   24*2048+ 696,   45*2048+ 697,   45*2048+ 698, 
  32*2048+ 702,    6*2048+ 703,   45*2048+ 704,   45*2048+ 705, 
  19*2048+ 706,   30*2048+ 707,   45*2048+ 708,   45*2048+ 709, 
   8*2048+ 710,   28*2048+ 711,   45*2048+ 712,   45*2048+ 713, 
   8*2048+ 714,   36*2048+ 715,   45*2048+ 716,   45*2048+ 717, 
  35*2048+ 718,   23*2048+ 719,   45*2048+ 720,   45*2048+ 721, 
  11*2048+ 722,   28*2048+ 723,   45*2048+ 724,   45*2048+ 725, 
  44*2048+ 735,   16*2048+ 736,   45*2048+ 737,   45*2048+ 738, 
   9*2048+ 739,    6*2048+ 740,   45*2048+ 741,   45*2048+ 742, 
   8*2048+ 743,    1*2048+ 744,   45*2048+ 745,   45*2048+ 746, 
  19*2048+ 747,   35*2048+ 748,   45*2048+ 749,   45*2048+ 750, 
  33*2048+ 754,    9*2048+ 755,   45*2048+ 756,   45*2048+ 757, 
   4*2048+ 758,   34*2048+ 759,   45*2048+ 760,   45*2048+ 761, 
  26*2048+ 762,   25*2048+ 763,   45*2048+ 764,   45*2048+ 765, 
  25*2048+ 766,   27*2048+ 767,   45*2048+ 768,   45*2048+ 769, 
   3*2048+ 770,    4*2048+ 771,   45*2048+ 772,   45*2048+ 773, 
  31*2048+ 783,    2*2048+ 784,   45*2048+ 785,   45*2048+ 786, 
  23*2048+ 790,   22*2048+ 791,   45*2048+ 792,   45*2048+ 793, 
   7*2048+ 794,   18*2048+ 795,   45*2048+ 796,   45*2048+ 797, 
  24*2048+ 798,   13*2048+ 799,   45*2048+ 800,   45*2048+ 801, 
  15*2048+ 802,    3*2048+ 803,   45*2048+ 804,   45*2048+ 805, 
   8*2048+ 806,   36*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  45*2048+ 810,   32*2048+ 811,   45*2048+ 812,   45*2048+ 813, 
  34*2048+ 814,   22*2048+ 815,   45*2048+ 816,   45*2048+ 817, 
   7*2048+ 818,   33*2048+ 819,   45*2048+ 820,   45*2048+ 821, 
  20*2048+ 822,   37*2048+ 823,   45*2048+ 824,   45*2048+ 825, 
  40*2048+ 826,   28*2048+ 827,   45*2048+ 828,   45*2048+ 829, 
  25*2048+ 830,   17*2048+ 831,   45*2048+ 832,   45*2048+ 833, 
  32*2048+ 837,    6*2048+ 838,   45*2048+ 839,   45*2048+ 840, 
  19*2048+ 841,   30*2048+ 842,   45*2048+ 843,   45*2048+ 844, 
   8*2048+ 845,   28*2048+ 846,   45*2048+ 847,   45*2048+ 848, 
   8*2048+ 849,   36*2048+ 850,   45*2048+ 851,   45*2048+ 852, 
  35*2048+ 853,   23*2048+ 854,   45*2048+ 855,   45*2048+ 856, 
  11*2048+ 857,   28*2048+ 858,   45*2048+ 859,   45*2048+ 860, 
  17*2048+ 870,   44*2048+ 871,   45*2048+ 872,   45*2048+ 873, 
  10*2048+ 874,    7*2048+ 875,   45*2048+ 876,   45*2048+ 877, 
   8*2048+ 878,    1*2048+ 879,   45*2048+ 880,   45*2048+ 881, 
  19*2048+ 882,   35*2048+ 883,   45*2048+ 884,   45*2048+ 885, 
  33*2048+ 889,    9*2048+ 890,   45*2048+ 891,   45*2048+ 892, 
   4*2048+ 893,   34*2048+ 894,   45*2048+ 895,   45*2048+ 896, 
  26*2048+ 897,   25*2048+ 898,   45*2048+ 899,   45*2048+ 900, 
  25*2048+ 901,   27*2048+ 902,   45*2048+ 903,   45*2048+ 904, 
   3*2048+ 905,    4*2048+ 906,   45*2048+ 907,   45*2048+ 908, 
  31*2048+ 918,    2*2048+ 919,   45*2048+ 920,   45*2048+ 921, 
  24*2048+ 925,   23*2048+ 926,   45*2048+ 927,   45*2048+ 928, 
   7*2048+ 929,   18*2048+ 930,   45*2048+ 931,   45*2048+ 932, 
  24*2048+ 933,   13*2048+ 934,   45*2048+ 935,   45*2048+ 936, 
  15*2048+ 937,    3*2048+ 938,   45*2048+ 939,   45*2048+ 940, 
   8*2048+ 941,   36*2048+ 942,   45*2048+ 943,   45*2048+ 944, 
  33*2048+ 945,   45*2048+ 946,   45*2048+ 947,   45*2048+ 948, 
  34*2048+ 949,   22*2048+ 950,   45*2048+ 951,   45*2048+ 952, 
   7*2048+ 953,   33*2048+ 954,   45*2048+ 955,   45*2048+ 956, 
  20*2048+ 957,   37*2048+ 958,   45*2048+ 959,   45*2048+ 960, 
  40*2048+ 961,   28*2048+ 962,   45*2048+ 963,   45*2048+ 964, 
  25*2048+ 965,   17*2048+ 966,   45*2048+ 967,   45*2048+ 968, 
   7*2048+ 972,   32*2048+ 973,   45*2048+ 974,   45*2048+ 975, 
  31*2048+ 976,   19*2048+ 977,   45*2048+ 978,   45*2048+ 979, 
   8*2048+ 980,   28*2048+ 981,   45*2048+ 982,   45*2048+ 983, 
   8*2048+ 984,   36*2048+ 985,   45*2048+ 986,   45*2048+ 987, 
  35*2048+ 988,   23*2048+ 989,   45*2048+ 990,   45*2048+ 991, 
  11*2048+ 992,   28*2048+ 993,   45*2048+ 994,   45*2048+ 995, 
  17*2048+1005,   44*2048+1006,   45*2048+1007,   45*2048+1008, 
  10*2048+1009,    7*2048+1010,   45*2048+1011,   45*2048+1012, 
   8*2048+1013,    1*2048+1014,   45*2048+1015,   45*2048+1016, 
  19*2048+1017,   35*2048+1018,   45*2048+1019,   45*2048+1020, 
  33*2048+1024,    9*2048+1025,   45*2048+1026,   45*2048+1027, 
   4*2048+1028,   34*2048+1029,   45*2048+1030,   45*2048+1031, 
  26*2048+1032,   26*2048+1033,   45*2048+1034,   45*2048+1035, 
  25*2048+1036,   27*2048+1037,   45*2048+1038,   45*2048+1039, 
   3*2048+1040,    4*2048+1041,   45*2048+1042,   45*2048+1043, 
  31*2048+1053,    2*2048+1054,   45*2048+1055,   45*2048+1056, 
  24*2048+1060,   23*2048+1061,   45*2048+1062,   45*2048+1063, 
   7*2048+1064,   18*2048+1065,   45*2048+1066,   45*2048+1067, 
  24*2048+1068,   13*2048+1069,   45*2048+1070,   45*2048+1071, 
  15*2048+1072,    3*2048+1073,   45*2048+1074,   45*2048+1075, 
   8*2048+1076,   36*2048+1077,   45*2048+1078,   45*2048+1079, 

  29*2048+   0,   27*2048+   1,    3*2048+   2,   45*2048+   3,   44*2048+   4, 
   9*2048+   5,   37*2048+   6,   19*2048+   7,   45*2048+   8,   45*2048+   9, 
  15*2048+  10,    1*2048+  11,   32*2048+  12,   45*2048+  13,   45*2048+  14, 
  17*2048+  15,   13*2048+  16,   29*2048+  17,   45*2048+  18,   45*2048+  19, 
  31*2048+  20,   40*2048+  21,   37*2048+  22,   45*2048+  23,   45*2048+  24, 
  30*2048+  25,   19*2048+  26,   38*2048+  27,   45*2048+  28,   45*2048+  29, 
  18*2048+  30,   31*2048+  31,   35*2048+  32,   45*2048+  33,   45*2048+  34, 
  33*2048+  35,    2*2048+  36,   33*2048+  37,   45*2048+  38,   45*2048+  39, 
   7*2048+  40,   12*2048+  41,   28*2048+  42,   45*2048+  43,   45*2048+  44, 
   5*2048+  45,    3*2048+  46,   23*2048+  47,   45*2048+  48,   45*2048+  49, 
   2*2048+  50,   34*2048+  51,   23*2048+  52,   45*2048+  53,   45*2048+  54, 
  32*2048+  55,   35*2048+  56,   28*2048+  57,   45*2048+  58,   45*2048+  59, 
  16*2048+  60,    6*2048+  61,   21*2048+  62,   45*2048+  63,   45*2048+  64, 
   9*2048+  65,   16*2048+  66,   22*2048+  67,   45*2048+  68,   45*2048+  69, 
  43*2048+  70,   41*2048+  71,   24*2048+  72,   45*2048+  73,   45*2048+  74, 
  18*2048+  75,   38*2048+  76,   36*2048+  77,   45*2048+  78,   45*2048+  79, 
  27*2048+  80,   27*2048+  81,    8*2048+  82,   45*2048+  83,   45*2048+  84, 
  10*2048+  85,   32*2048+  86,    2*2048+  87,   45*2048+  88,   45*2048+  89, 
  24*2048+  90,    3*2048+  91,    2*2048+  92,   45*2048+  93,   45*2048+  94, 
  27*2048+  95,   24*2048+  96,   24*2048+  97,   45*2048+  98,   45*2048+  99, 
  22*2048+ 100,   19*2048+ 101,   16*2048+ 102,   45*2048+ 103,   45*2048+ 104, 
  37*2048+ 105,   30*2048+ 106,   14*2048+ 107,   45*2048+ 108,   45*2048+ 109, 
  26*2048+ 110,   30*2048+ 111,   32*2048+ 112,   45*2048+ 113,   45*2048+ 114, 
  31*2048+ 115,   42*2048+ 116,   17*2048+ 117,   45*2048+ 118,   45*2048+ 119, 
   6*2048+ 120,   26*2048+ 121,   14*2048+ 122,   45*2048+ 123,   45*2048+ 124, 
  22*2048+ 125,   13*2048+ 126,   30*2048+ 127,   45*2048+ 128,   45*2048+ 129, 
  43*2048+ 130,   30*2048+ 131,   24*2048+ 132,   45*2048+ 133,   45*2048+ 134, 
   3*2048+ 135,   15*2048+ 136,   31*2048+ 137,   45*2048+ 138,   45*2048+ 139, 
   6*2048+ 140,   25*2048+ 141,   14*2048+ 142,   45*2048+ 143,   45*2048+ 144, 
   8*2048+ 145,    9*2048+ 146,    5*2048+ 147,   45*2048+ 148,   45*2048+ 149, 
  29*2048+ 150,   27*2048+ 151,    3*2048+ 152,   45*2048+ 153,   45*2048+ 154, 
  20*2048+ 155,    9*2048+ 156,   37*2048+ 157,   45*2048+ 158,   45*2048+ 159, 
  33*2048+ 160,   15*2048+ 161,    1*2048+ 162,   45*2048+ 163,   45*2048+ 164, 
  17*2048+ 165,   13*2048+ 166,   29*2048+ 167,   45*2048+ 168,   45*2048+ 169, 
  38*2048+ 170,   31*2048+ 171,   40*2048+ 172,   45*2048+ 173,   45*2048+ 174, 
  30*2048+ 175,   19*2048+ 176,   38*2048+ 177,   45*2048+ 178,   45*2048+ 179, 
  18*2048+ 180,   31*2048+ 181,   35*2048+ 182,   45*2048+ 183,   45*2048+ 184, 
  33*2048+ 185,    2*2048+ 186,   33*2048+ 187,   45*2048+ 188,   45*2048+ 189, 
  29*2048+ 190,    7*2048+ 191,   12*2048+ 192,   45*2048+ 193,   45*2048+ 194, 
   5*2048+ 195,    3*2048+ 196,   23*2048+ 197,   45*2048+ 198,   45*2048+ 199, 
   2*2048+ 200,   34*2048+ 201,   23*2048+ 202,   45*2048+ 203,   45*2048+ 204, 
  32*2048+ 205,   35*2048+ 206,   28*2048+ 207,   45*2048+ 208,   45*2048+ 209, 
  16*2048+ 210,    6*2048+ 211,   21*2048+ 212,   45*2048+ 213,   45*2048+ 214, 
   9*2048+ 215,   16*2048+ 216,   22*2048+ 217,   45*2048+ 218,   45*2048+ 219, 
  25*2048+ 220,   43*2048+ 221,   41*2048+ 222,   45*2048+ 223,   45*2048+ 224, 
  37*2048+ 225,   18*2048+ 226,   38*2048+ 227,   45*2048+ 228,   45*2048+ 229, 
  27*2048+ 230,   27*2048+ 231,    8*2048+ 232,   45*2048+ 233,   45*2048+ 234, 
   3*2048+ 235,   10*2048+ 236,   32*2048+ 237,   45*2048+ 238,   45*2048+ 239, 
  24*2048+ 240,    3*2048+ 241,    2*2048+ 242,   45*2048+ 243,   45*2048+ 244, 
  27*2048+ 245,   24*2048+ 246,   24*2048+ 247,   45*2048+ 248,   45*2048+ 249, 
  22*2048+ 250,   19*2048+ 251,   16*2048+ 252,   45*2048+ 253,   45*2048+ 254, 
  37*2048+ 255,   30*2048+ 256,   14*2048+ 257,   45*2048+ 258,   45*2048+ 259, 
  26*2048+ 260,   30*2048+ 261,   32*2048+ 262,   45*2048+ 263,   45*2048+ 264, 
  31*2048+ 265,   42*2048+ 266,   17*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
   6*2048+ 270,   26*2048+ 271,   14*2048+ 272,   45*2048+ 273,   45*2048+ 274, 
  22*2048+ 275,   13*2048+ 276,   30*2048+ 277,   45*2048+ 278,   45*2048+ 279, 
  43*2048+ 280,   30*2048+ 281,   24*2048+ 282,   45*2048+ 283,   45*2048+ 284, 
   3*2048+ 285,   15*2048+ 286,   31*2048+ 287,   45*2048+ 288,   45*2048+ 289, 
   6*2048+ 290,   25*2048+ 291,   14*2048+ 292,   45*2048+ 293,   45*2048+ 294, 
   8*2048+ 295,    9*2048+ 296,    5*2048+ 297,   45*2048+ 298,   45*2048+ 299, 
  29*2048+ 300,   27*2048+ 301,    3*2048+ 302,   45*2048+ 303,   45*2048+ 304, 
  20*2048+ 305,    9*2048+ 306,   37*2048+ 307,   45*2048+ 308,   45*2048+ 309, 
  33*2048+ 310,   15*2048+ 311,    1*2048+ 312,   45*2048+ 313,   45*2048+ 314, 
  17*2048+ 315,   13*2048+ 316,   29*2048+ 317,   45*2048+ 318,   45*2048+ 319, 
  38*2048+ 320,   31*2048+ 321,   40*2048+ 322,   45*2048+ 323,   45*2048+ 324, 
  39*2048+ 325,   30*2048+ 326,   19*2048+ 327,   45*2048+ 328,   45*2048+ 329, 
  36*2048+ 330,   18*2048+ 331,   31*2048+ 332,   45*2048+ 333,   45*2048+ 334, 
   3*2048+ 335,   34*2048+ 336,   33*2048+ 337,   45*2048+ 338,   45*2048+ 339, 
  29*2048+ 340,    7*2048+ 341,   12*2048+ 342,   45*2048+ 343,   45*2048+ 344, 
   5*2048+ 345,    3*2048+ 346,   23*2048+ 347,   45*2048+ 348,   45*2048+ 349, 
   2*2048+ 350,   34*2048+ 351,   23*2048+ 352,   45*2048+ 353,   45*2048+ 354, 
  32*2048+ 355,   35*2048+ 356,   28*2048+ 357,   45*2048+ 358,   45*2048+ 359, 
  16*2048+ 360,    6*2048+ 361,   21*2048+ 362,   45*2048+ 363,   45*2048+ 364, 
   9*2048+ 365,   16*2048+ 366,   22*2048+ 367,   45*2048+ 368,   45*2048+ 369, 
  25*2048+ 370,   43*2048+ 371,   41*2048+ 372,   45*2048+ 373,   45*2048+ 374, 
  39*2048+ 375,   37*2048+ 376,   18*2048+ 377,   45*2048+ 378,   45*2048+ 379, 
  28*2048+ 380,    9*2048+ 381,   27*2048+ 382,   45*2048+ 383,   45*2048+ 384, 
  33*2048+ 385,    3*2048+ 386,   10*2048+ 387,   45*2048+ 388,   45*2048+ 389, 
  24*2048+ 390,    3*2048+ 391,    2*2048+ 392,   45*2048+ 393,   45*2048+ 394, 
  25*2048+ 395,   27*2048+ 396,   24*2048+ 397,   45*2048+ 398,   45*2048+ 399, 
  22*2048+ 400,   19*2048+ 401,   16*2048+ 402,   45*2048+ 403,   45*2048+ 404, 
  31*2048+ 405,   15*2048+ 406,   37*2048+ 407,   45*2048+ 408,   45*2048+ 409, 
  26*2048+ 410,   30*2048+ 411,   32*2048+ 412,   45*2048+ 413,   45*2048+ 414, 
  31*2048+ 415,   42*2048+ 416,   17*2048+ 417,   45*2048+ 418,   45*2048+ 419, 
   6*2048+ 420,   26*2048+ 421,   14*2048+ 422,   45*2048+ 423,   45*2048+ 424, 
  22*2048+ 425,   13*2048+ 426,   30*2048+ 427,   45*2048+ 428,   45*2048+ 429, 
  43*2048+ 430,   30*2048+ 431,   24*2048+ 432,   45*2048+ 433,   45*2048+ 434, 
   3*2048+ 435,   15*2048+ 436,   31*2048+ 437,   45*2048+ 438,   45*2048+ 439, 
  15*2048+ 440,    6*2048+ 441,   25*2048+ 442,   45*2048+ 443,   45*2048+ 444, 
   8*2048+ 445,    9*2048+ 446,    5*2048+ 447,   45*2048+ 448,   45*2048+ 449, 
   4*2048+ 450,   29*2048+ 451,   27*2048+ 452,   45*2048+ 453,   45*2048+ 454, 
  20*2048+ 455,    9*2048+ 456,   37*2048+ 457,   45*2048+ 458,   45*2048+ 459, 
  33*2048+ 460,   15*2048+ 461,    1*2048+ 462,   45*2048+ 463,   45*2048+ 464, 
  30*2048+ 465,   17*2048+ 466,   13*2048+ 467,   45*2048+ 468,   45*2048+ 469, 
  38*2048+ 470,   31*2048+ 471,   40*2048+ 472,   45*2048+ 473,   45*2048+ 474, 
  39*2048+ 475,   30*2048+ 476,   19*2048+ 477,   45*2048+ 478,   45*2048+ 479, 
  32*2048+ 480,   36*2048+ 481,   18*2048+ 482,   45*2048+ 483,   45*2048+ 484, 
   3*2048+ 485,   34*2048+ 486,   33*2048+ 487,   45*2048+ 488,   45*2048+ 489, 
   8*2048+ 490,   13*2048+ 491,   29*2048+ 492,   45*2048+ 493,   45*2048+ 494, 
  24*2048+ 495,    5*2048+ 496,    3*2048+ 497,   45*2048+ 498,   45*2048+ 499, 
  24*2048+ 500,    2*2048+ 501,   34*2048+ 502,   45*2048+ 503,   45*2048+ 504, 
  29*2048+ 505,   32*2048+ 506,   35*2048+ 507,   45*2048+ 508,   45*2048+ 509, 
  16*2048+ 510,    6*2048+ 511,   21*2048+ 512,   45*2048+ 513,   45*2048+ 514, 
  23*2048+ 515,    9*2048+ 516,   16*2048+ 517,   45*2048+ 518,   45*2048+ 519, 
  25*2048+ 520,   43*2048+ 521,   41*2048+ 522,   45*2048+ 523,   45*2048+ 524, 
  39*2048+ 525,   37*2048+ 526,   18*2048+ 527,   45*2048+ 528,   45*2048+ 529, 
  28*2048+ 530,    9*2048+ 531,   27*2048+ 532,   45*2048+ 533,   45*2048+ 534, 
  11*2048+ 535,   33*2048+ 536,    3*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
  24*2048+ 540,    3*2048+ 541,    2*2048+ 542,   45*2048+ 543,   45*2048+ 544, 
  25*2048+ 545,   27*2048+ 546,   24*2048+ 547,   45*2048+ 548,   45*2048+ 549, 
  20*2048+ 550,   17*2048+ 551,   22*2048+ 552,   45*2048+ 553,   45*2048+ 554, 
  31*2048+ 555,   15*2048+ 556,   37*2048+ 557,   45*2048+ 558,   45*2048+ 559, 
  26*2048+ 560,   30*2048+ 561,   32*2048+ 562,   45*2048+ 563,   45*2048+ 564, 
  31*2048+ 565,   42*2048+ 566,   17*2048+ 567,   45*2048+ 568,   45*2048+ 569, 
   6*2048+ 570,   26*2048+ 571,   14*2048+ 572,   45*2048+ 573,   45*2048+ 574, 
  22*2048+ 575,   13*2048+ 576,   30*2048+ 577,   45*2048+ 578,   45*2048+ 579, 
  43*2048+ 580,   30*2048+ 581,   24*2048+ 582,   45*2048+ 583,   45*2048+ 584, 
  16*2048+ 585,   32*2048+ 586,    3*2048+ 587,   45*2048+ 588,   45*2048+ 589, 
  15*2048+ 590,    6*2048+ 591,   25*2048+ 592,   45*2048+ 593,   45*2048+ 594, 
   8*2048+ 595,    9*2048+ 596,    5*2048+ 597,   45*2048+ 598,   45*2048+ 599, 
   4*2048+ 600,   29*2048+ 601,   27*2048+ 602,   45*2048+ 603,   45*2048+ 604, 
  20*2048+ 605,    9*2048+ 606,   37*2048+ 607,   45*2048+ 608,   45*2048+ 609, 
  33*2048+ 610,   15*2048+ 611,    1*2048+ 612,   45*2048+ 613,   45*2048+ 614, 
  14*2048+ 615,   30*2048+ 616,   17*2048+ 617,   45*2048+ 618,   45*2048+ 619, 
  38*2048+ 620,   31*2048+ 621,   40*2048+ 622,   45*2048+ 623,   45*2048+ 624, 
  39*2048+ 625,   30*2048+ 626,   19*2048+ 627,   45*2048+ 628,   45*2048+ 629, 
  32*2048+ 630,   36*2048+ 631,   18*2048+ 632,   45*2048+ 633,   45*2048+ 634, 
   3*2048+ 635,   34*2048+ 636,   33*2048+ 637,   45*2048+ 638,   45*2048+ 639, 
   8*2048+ 640,   13*2048+ 641,   29*2048+ 642,   45*2048+ 643,   45*2048+ 644, 
  24*2048+ 645,    5*2048+ 646,    3*2048+ 647,   45*2048+ 648,   45*2048+ 649, 
  24*2048+ 650,    2*2048+ 651,   34*2048+ 652,   45*2048+ 653,   45*2048+ 654, 
  33*2048+ 655,   36*2048+ 656,   29*2048+ 657,   45*2048+ 658,   45*2048+ 659, 
  16*2048+ 660,    6*2048+ 661,   21*2048+ 662,   45*2048+ 663,   45*2048+ 664, 
  23*2048+ 665,    9*2048+ 666,   16*2048+ 667,   45*2048+ 668,   45*2048+ 669, 
  25*2048+ 670,   43*2048+ 671,   41*2048+ 672,   45*2048+ 673,   45*2048+ 674, 
  39*2048+ 675,   37*2048+ 676,   18*2048+ 677,   45*2048+ 678,   45*2048+ 679, 
  28*2048+ 680,    9*2048+ 681,   27*2048+ 682,   45*2048+ 683,   45*2048+ 684, 
  11*2048+ 685,   33*2048+ 686,    3*2048+ 687,   45*2048+ 688,   45*2048+ 689, 
   3*2048+ 690,   24*2048+ 691,    3*2048+ 692,   45*2048+ 693,   45*2048+ 694, 
  25*2048+ 695,   27*2048+ 696,   24*2048+ 697,   45*2048+ 698,   45*2048+ 699, 
  23*2048+ 700,   20*2048+ 701,   17*2048+ 702,   45*2048+ 703,   45*2048+ 704, 
  31*2048+ 705,   15*2048+ 706,   37*2048+ 707,   45*2048+ 708,   45*2048+ 709, 
  26*2048+ 710,   30*2048+ 711,   32*2048+ 712,   45*2048+ 713,   45*2048+ 714, 
  18*2048+ 715,   31*2048+ 716,   42*2048+ 717,   45*2048+ 718,   45*2048+ 719, 
   6*2048+ 720,   26*2048+ 721,   14*2048+ 722,   45*2048+ 723,   45*2048+ 724, 
  31*2048+ 725,   22*2048+ 726,   13*2048+ 727,   45*2048+ 728,   45*2048+ 729, 
  25*2048+ 730,   43*2048+ 731,   30*2048+ 732,   45*2048+ 733,   45*2048+ 734, 
  16*2048+ 735,   32*2048+ 736,    3*2048+ 737,   45*2048+ 738,   45*2048+ 739, 
  15*2048+ 740,    6*2048+ 741,   25*2048+ 742,   45*2048+ 743,   45*2048+ 744, 
   8*2048+ 745,    9*2048+ 746,    5*2048+ 747,   45*2048+ 748,   45*2048+ 749, 
   4*2048+ 750,   29*2048+ 751,   27*2048+ 752,   45*2048+ 753,   45*2048+ 754, 
  10*2048+ 755,   38*2048+ 756,   20*2048+ 757,   45*2048+ 758,   45*2048+ 759, 
   2*2048+ 760,   33*2048+ 761,   15*2048+ 762,   45*2048+ 763,   45*2048+ 764, 
  14*2048+ 765,   30*2048+ 766,   17*2048+ 767,   45*2048+ 768,   45*2048+ 769, 
  41*2048+ 770,   38*2048+ 771,   31*2048+ 772,   45*2048+ 773,   45*2048+ 774, 
  39*2048+ 775,   30*2048+ 776,   19*2048+ 777,   45*2048+ 778,   45*2048+ 779, 
  19*2048+ 780,   32*2048+ 781,   36*2048+ 782,   45*2048+ 783,   45*2048+ 784, 
  34*2048+ 785,    3*2048+ 786,   34*2048+ 787,   45*2048+ 788,   45*2048+ 789, 
   8*2048+ 790,   13*2048+ 791,   29*2048+ 792,   45*2048+ 793,   45*2048+ 794, 
  24*2048+ 795,    5*2048+ 796,    3*2048+ 797,   45*2048+ 798,   45*2048+ 799, 
  35*2048+ 800,   24*2048+ 801,    2*2048+ 802,   45*2048+ 803,   45*2048+ 804, 
  33*2048+ 805,   36*2048+ 806,   29*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  22*2048+ 810,   16*2048+ 811,    6*2048+ 812,   45*2048+ 813,   45*2048+ 814, 
  17*2048+ 815,   23*2048+ 816,    9*2048+ 817,   45*2048+ 818,   45*2048+ 819, 
  25*2048+ 820,   43*2048+ 821,   41*2048+ 822,   45*2048+ 823,   45*2048+ 824, 
  19*2048+ 825,   39*2048+ 826,   37*2048+ 827,   45*2048+ 828,   45*2048+ 829, 
  28*2048+ 830,    9*2048+ 831,   27*2048+ 832,   45*2048+ 833,   45*2048+ 834, 
  11*2048+ 835,   33*2048+ 836,    3*2048+ 837,   45*2048+ 838,   45*2048+ 839, 
   4*2048+ 840,    3*2048+ 841,   24*2048+ 842,   45*2048+ 843,   45*2048+ 844, 
  25*2048+ 845,   25*2048+ 846,   27*2048+ 847,   45*2048+ 848,   45*2048+ 849, 
  23*2048+ 850,   20*2048+ 851,   17*2048+ 852,   45*2048+ 853,   45*2048+ 854, 
  31*2048+ 855,   15*2048+ 856,   37*2048+ 857,   45*2048+ 858,   45*2048+ 859, 
  26*2048+ 860,   30*2048+ 861,   32*2048+ 862,   45*2048+ 863,   45*2048+ 864, 
  18*2048+ 865,   31*2048+ 866,   42*2048+ 867,   45*2048+ 868,   45*2048+ 869, 
   6*2048+ 870,   26*2048+ 871,   14*2048+ 872,   45*2048+ 873,   45*2048+ 874, 
  14*2048+ 875,   31*2048+ 876,   22*2048+ 877,   45*2048+ 878,   45*2048+ 879, 
  44*2048+ 880,   31*2048+ 881,   25*2048+ 882,   45*2048+ 883,   45*2048+ 884, 
   4*2048+ 885,   16*2048+ 886,   32*2048+ 887,   45*2048+ 888,   45*2048+ 889, 
  15*2048+ 890,    6*2048+ 891,   25*2048+ 892,   45*2048+ 893,   45*2048+ 894, 
   8*2048+ 895,    9*2048+ 896,    5*2048+ 897,   45*2048+ 898,   45*2048+ 899, 
   4*2048+ 900,   29*2048+ 901,   27*2048+ 902,   45*2048+ 903,   45*2048+ 904, 
  10*2048+ 905,   38*2048+ 906,   20*2048+ 907,   45*2048+ 908,   45*2048+ 909, 
   2*2048+ 910,   33*2048+ 911,   15*2048+ 912,   45*2048+ 913,   45*2048+ 914, 
  14*2048+ 915,   30*2048+ 916,   17*2048+ 917,   45*2048+ 918,   45*2048+ 919, 
  41*2048+ 920,   38*2048+ 921,   31*2048+ 922,   45*2048+ 923,   45*2048+ 924, 
  39*2048+ 925,   30*2048+ 926,   19*2048+ 927,   45*2048+ 928,   45*2048+ 929, 
  19*2048+ 930,   32*2048+ 931,   36*2048+ 932,   45*2048+ 933,   45*2048+ 934, 
  34*2048+ 935,    3*2048+ 936,   34*2048+ 937,   45*2048+ 938,   45*2048+ 939, 
   8*2048+ 940,   13*2048+ 941,   29*2048+ 942,   45*2048+ 943,   45*2048+ 944, 
  24*2048+ 945,    5*2048+ 946,    3*2048+ 947,   45*2048+ 948,   45*2048+ 949, 
   3*2048+ 950,   35*2048+ 951,   24*2048+ 952,   45*2048+ 953,   45*2048+ 954, 
  33*2048+ 955,   36*2048+ 956,   29*2048+ 957,   45*2048+ 958,   45*2048+ 959, 
  17*2048+ 960,    7*2048+ 961,   22*2048+ 962,   45*2048+ 963,   45*2048+ 964, 
  10*2048+ 965,   17*2048+ 966,   23*2048+ 967,   45*2048+ 968,   45*2048+ 969, 
  44*2048+ 970,   42*2048+ 971,   25*2048+ 972,   45*2048+ 973,   45*2048+ 974, 
  19*2048+ 975,   39*2048+ 976,   37*2048+ 977,   45*2048+ 978,   45*2048+ 979, 
  28*2048+ 980,    9*2048+ 981,   27*2048+ 982,   45*2048+ 983,   45*2048+ 984, 
  11*2048+ 985,   33*2048+ 986,    3*2048+ 987,   45*2048+ 988,   45*2048+ 989, 
   4*2048+ 990,    3*2048+ 991,   24*2048+ 992,   45*2048+ 993,   45*2048+ 994, 
  25*2048+ 995,   25*2048+ 996,   27*2048+ 997,   45*2048+ 998,   45*2048+ 999, 
  23*2048+1000,   20*2048+1001,   17*2048+1002,   45*2048+1003,   45*2048+1004, 
  31*2048+1005,   15*2048+1006,   37*2048+1007,   45*2048+1008,   45*2048+1009, 
  26*2048+1010,   30*2048+1011,   32*2048+1012,   45*2048+1013,   45*2048+1014, 
  18*2048+1015,   31*2048+1016,   42*2048+1017,   45*2048+1018,   45*2048+1019, 
  15*2048+1020,    6*2048+1021,   26*2048+1022,   45*2048+1023,   45*2048+1024, 
  23*2048+1025,   14*2048+1026,   31*2048+1027,   45*2048+1028,   45*2048+1029, 
  44*2048+1030,   31*2048+1031,   25*2048+1032,   45*2048+1033,   45*2048+1034, 
   4*2048+1035,   16*2048+1036,   32*2048+1037,   45*2048+1038,   45*2048+1039, 
  26*2048+1040,   15*2048+1041,    6*2048+1042,   45*2048+1043,   45*2048+1044, 
   6*2048+1045,    8*2048+1046,    9*2048+1047,   45*2048+1048,   45*2048+1049, 
  28*2048+1050,    4*2048+1051,   29*2048+1052,   45*2048+1053,   45*2048+1054, 
  10*2048+1055,   38*2048+1056,   20*2048+1057,   45*2048+1058,   45*2048+1059, 
  16*2048+1060,    2*2048+1061,   33*2048+1062,   45*2048+1063,   45*2048+1064, 
  14*2048+1065,   30*2048+1066,   17*2048+1067,   45*2048+1068,   45*2048+1069, 
  32*2048+1070,   41*2048+1071,   38*2048+1072,   45*2048+1073,   45*2048+1074, 
  31*2048+1075,   20*2048+1076,   39*2048+1077,   45*2048+1078,   45*2048+1079, 
  19*2048+1080,   32*2048+1081,   36*2048+1082,   45*2048+1083,   45*2048+1084, 
  34*2048+1085,    3*2048+1086,   34*2048+1087,   45*2048+1088,   45*2048+1089, 
   8*2048+1090,   13*2048+1091,   29*2048+1092,   45*2048+1093,   45*2048+1094, 
   4*2048+1095,   24*2048+1096,    5*2048+1097,   45*2048+1098,   45*2048+1099, 
   3*2048+1100,   35*2048+1101,   24*2048+1102,   45*2048+1103,   45*2048+1104, 
  33*2048+1105,   36*2048+1106,   29*2048+1107,   45*2048+1108,   45*2048+1109, 
  17*2048+1110,    7*2048+1111,   22*2048+1112,   45*2048+1113,   45*2048+1114, 
  10*2048+1115,   17*2048+1116,   23*2048+1117,   45*2048+1118,   45*2048+1119, 
  44*2048+1120,   42*2048+1121,   25*2048+1122,   45*2048+1123,   45*2048+1124, 
  19*2048+1125,   39*2048+1126,   37*2048+1127,   45*2048+1128,   45*2048+1129, 
  28*2048+1130,   28*2048+1131,    9*2048+1132,   45*2048+1133,   45*2048+1134, 
  11*2048+1135,   33*2048+1136,    3*2048+1137,   45*2048+1138,   45*2048+1139, 
   4*2048+1140,    3*2048+1141,   24*2048+1142,   45*2048+1143,   45*2048+1144, 
  25*2048+1145,   25*2048+1146,   27*2048+1147,   45*2048+1148,   45*2048+1149, 
  23*2048+1150,   20*2048+1151,   17*2048+1152,   45*2048+1153,   45*2048+1154, 
  31*2048+1155,   15*2048+1156,   37*2048+1157,   45*2048+1158,   45*2048+1159, 
  33*2048+1160,   26*2048+1161,   30*2048+1162,   45*2048+1163,   45*2048+1164, 
  18*2048+1165,   31*2048+1166,   42*2048+1167,   45*2048+1168,   45*2048+1169, 
  27*2048+1170,   15*2048+1171,    6*2048+1172,   45*2048+1173,   45*2048+1174, 
  23*2048+1175,   14*2048+1176,   31*2048+1177,   45*2048+1178,   45*2048+1179, 
  44*2048+1180,   31*2048+1181,   25*2048+1182,   45*2048+1183,   45*2048+1184, 
   4*2048+1185,   16*2048+1186,   32*2048+1187,   45*2048+1188,   45*2048+1189, 
  26*2048+1190,   15*2048+1191,    6*2048+1192,   45*2048+1193,   45*2048+1194, 
   6*2048+1195,    8*2048+1196,    9*2048+1197,   45*2048+1198,   45*2048+1199, 

   0*2048+   0,   24*2048+   1,   43*2048+   2,    3*2048+   3,   45*2048+   4,   44*2048+   5, 
  27*2048+   6,   23*2048+   7,   21*2048+   8,   13*2048+   9,   45*2048+  10,   45*2048+  11, 
  20*2048+  12,    4*2048+  13,   30*2048+  14,   36*2048+  15,   45*2048+  16,   45*2048+  17, 
  13*2048+  18,   36*2048+  19,   34*2048+  20,   18*2048+  21,   45*2048+  22,   45*2048+  23, 
  26*2048+  24,   38*2048+  25,   21*2048+  26,    5*2048+  27,   45*2048+  28,   45*2048+  29, 
  22*2048+  30,   37*2048+  31,    8*2048+  32,   17*2048+  33,   45*2048+  34,   45*2048+  35, 
  15*2048+  36,    3*2048+  37,   13*2048+  38,    2*2048+  39,   45*2048+  40,   45*2048+  41, 
  26*2048+  42,   18*2048+  43,    1*2048+  44,   10*2048+  45,   45*2048+  46,   45*2048+  47, 
  25*2048+  48,    3*2048+  49,   16*2048+  50,   17*2048+  51,   45*2048+  52,   45*2048+  53, 
  33*2048+  54,   14*2048+  55,   41*2048+  56,   14*2048+  57,   45*2048+  58,   45*2048+  59, 
  13*2048+  60,   43*2048+  61,   21*2048+  62,   38*2048+  63,   45*2048+  64,   45*2048+  65, 
  44*2048+  66,   36*2048+  67,   37*2048+  68,   24*2048+  69,   45*2048+  70,   45*2048+  71, 
   4*2048+  72,   18*2048+  73,   25*2048+  74,   36*2048+  75,   45*2048+  76,   45*2048+  77, 
  33*2048+  78,   27*2048+  79,   34*2048+  80,   34*2048+  81,   45*2048+  82,   45*2048+  83, 
  42*2048+  84,   36*2048+  85,   42*2048+  86,   32*2048+  87,   45*2048+  88,   45*2048+  89, 
   2*2048+  90,   41*2048+  91,   36*2048+  92,    1*2048+  93,   45*2048+  94,   45*2048+  95, 
   9*2048+  96,   14*2048+  97,   42*2048+  98,    4*2048+  99,   45*2048+ 100,   45*2048+ 101, 
  10*2048+ 102,    9*2048+ 103,    7*2048+ 104,   36*2048+ 105,   45*2048+ 106,   45*2048+ 107, 
   7*2048+ 108,   26*2048+ 109,   29*2048+ 110,   22*2048+ 111,   45*2048+ 112,   45*2048+ 113, 
  19*2048+ 114,    4*2048+ 115,    1*2048+ 116,   27*2048+ 117,   45*2048+ 118,   45*2048+ 119, 
  41*2048+ 120,   24*2048+ 121,   36*2048+ 122,   24*2048+ 123,   45*2048+ 124,   45*2048+ 125, 
  30*2048+ 126,    0*2048+ 127,   24*2048+ 128,   38*2048+ 129,   45*2048+ 130,   45*2048+ 131, 
  41*2048+ 132,   23*2048+ 133,   11*2048+ 134,   35*2048+ 135,   45*2048+ 136,   45*2048+ 137, 
  20*2048+ 138,   41*2048+ 139,   26*2048+ 140,    5*2048+ 141,   45*2048+ 142,   45*2048+ 143, 
  14*2048+ 144,    8*2048+ 145,   41*2048+ 146,    3*2048+ 147,   45*2048+ 148,   45*2048+ 149, 
   2*2048+ 150,   11*2048+ 151,    4*2048+ 152,    7*2048+ 153,   45*2048+ 154,   45*2048+ 155, 
  12*2048+ 156,    3*2048+ 157,   18*2048+ 158,   10*2048+ 159,   45*2048+ 160,   45*2048+ 161, 
   0*2048+ 162,   24*2048+ 163,   43*2048+ 164,    3*2048+ 165,   45*2048+ 166,   45*2048+ 167, 
  14*2048+ 168,   27*2048+ 169,   23*2048+ 170,   21*2048+ 171,   45*2048+ 172,   45*2048+ 173, 
  20*2048+ 174,    4*2048+ 175,   30*2048+ 176,   36*2048+ 177,   45*2048+ 178,   45*2048+ 179, 
  35*2048+ 180,   19*2048+ 181,   13*2048+ 182,   36*2048+ 183,   45*2048+ 184,   45*2048+ 185, 
  26*2048+ 186,   38*2048+ 187,   21*2048+ 188,    5*2048+ 189,   45*2048+ 190,   45*2048+ 191, 
  18*2048+ 192,   22*2048+ 193,   37*2048+ 194,    8*2048+ 195,   45*2048+ 196,   45*2048+ 197, 
  15*2048+ 198,    3*2048+ 199,   13*2048+ 200,    2*2048+ 201,   45*2048+ 202,   45*2048+ 203, 
  19*2048+ 204,    2*2048+ 205,   11*2048+ 206,   26*2048+ 207,   45*2048+ 208,   45*2048+ 209, 
  18*2048+ 210,   25*2048+ 211,    3*2048+ 212,   16*2048+ 213,   45*2048+ 214,   45*2048+ 215, 
  33*2048+ 216,   14*2048+ 217,   41*2048+ 218,   14*2048+ 219,   45*2048+ 220,   45*2048+ 221, 
  13*2048+ 222,   43*2048+ 223,   21*2048+ 224,   38*2048+ 225,   45*2048+ 226,   45*2048+ 227, 
  44*2048+ 228,   36*2048+ 229,   37*2048+ 230,   24*2048+ 231,   45*2048+ 232,   45*2048+ 233, 
  26*2048+ 234,   37*2048+ 235,    4*2048+ 236,   18*2048+ 237,   45*2048+ 238,   45*2048+ 239, 
  33*2048+ 240,   27*2048+ 241,   34*2048+ 242,   34*2048+ 243,   45*2048+ 244,   45*2048+ 245, 
  42*2048+ 246,   36*2048+ 247,   42*2048+ 248,   32*2048+ 249,   45*2048+ 250,   45*2048+ 251, 
  37*2048+ 252,    2*2048+ 253,    2*2048+ 254,   41*2048+ 255,   45*2048+ 256,   45*2048+ 257, 
   5*2048+ 258,    9*2048+ 259,   14*2048+ 260,   42*2048+ 261,   45*2048+ 262,   45*2048+ 263, 
  10*2048+ 264,    9*2048+ 265,    7*2048+ 266,   36*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
   7*2048+ 270,   26*2048+ 271,   29*2048+ 272,   22*2048+ 273,   45*2048+ 274,   45*2048+ 275, 
  19*2048+ 276,    4*2048+ 277,    1*2048+ 278,   27*2048+ 279,   45*2048+ 280,   45*2048+ 281, 
  25*2048+ 282,   41*2048+ 283,   24*2048+ 284,   36*2048+ 285,   45*2048+ 286,   45*2048+ 287, 
  39*2048+ 288,   30*2048+ 289,    0*2048+ 290,   24*2048+ 291,   45*2048+ 292,   45*2048+ 293, 
  36*2048+ 294,   41*2048+ 295,   23*2048+ 296,   11*2048+ 297,   45*2048+ 298,   45*2048+ 299, 
   6*2048+ 300,   20*2048+ 301,   41*2048+ 302,   26*2048+ 303,   45*2048+ 304,   45*2048+ 305, 
  14*2048+ 306,    8*2048+ 307,   41*2048+ 308,    3*2048+ 309,   45*2048+ 310,   45*2048+ 311, 
   2*2048+ 312,   11*2048+ 313,    4*2048+ 314,    7*2048+ 315,   45*2048+ 316,   45*2048+ 317, 
  11*2048+ 318,   12*2048+ 319,    3*2048+ 320,   18*2048+ 321,   45*2048+ 322,   45*2048+ 323, 
   4*2048+ 324,    0*2048+ 325,   24*2048+ 326,   43*2048+ 327,   45*2048+ 328,   45*2048+ 329, 
  22*2048+ 330,   14*2048+ 331,   27*2048+ 332,   23*2048+ 333,   45*2048+ 334,   45*2048+ 335, 
  20*2048+ 336,    4*2048+ 337,   30*2048+ 338,   36*2048+ 339,   45*2048+ 340,   45*2048+ 341, 
  35*2048+ 342,   19*2048+ 343,   13*2048+ 344,   36*2048+ 345,   45*2048+ 346,   45*2048+ 347, 
  26*2048+ 348,   38*2048+ 349,   21*2048+ 350,    5*2048+ 351,   45*2048+ 352,   45*2048+ 353, 
  18*2048+ 354,   22*2048+ 355,   37*2048+ 356,    8*2048+ 357,   45*2048+ 358,   45*2048+ 359, 
  15*2048+ 360,    3*2048+ 361,   13*2048+ 362,    2*2048+ 363,   45*2048+ 364,   45*2048+ 365, 
  19*2048+ 366,    2*2048+ 367,   11*2048+ 368,   26*2048+ 369,   45*2048+ 370,   45*2048+ 371, 
  18*2048+ 372,   25*2048+ 373,    3*2048+ 374,   16*2048+ 375,   45*2048+ 376,   45*2048+ 377, 
  15*2048+ 378,   33*2048+ 379,   14*2048+ 380,   41*2048+ 381,   45*2048+ 382,   45*2048+ 383, 
  13*2048+ 384,   43*2048+ 385,   21*2048+ 386,   38*2048+ 387,   45*2048+ 388,   45*2048+ 389, 
  44*2048+ 390,   36*2048+ 391,   37*2048+ 392,   24*2048+ 393,   45*2048+ 394,   45*2048+ 395, 
  26*2048+ 396,   37*2048+ 397,    4*2048+ 398,   18*2048+ 399,   45*2048+ 400,   45*2048+ 401, 
  35*2048+ 402,   33*2048+ 403,   27*2048+ 404,   34*2048+ 405,   45*2048+ 406,   45*2048+ 407, 
  43*2048+ 408,   33*2048+ 409,   42*2048+ 410,   36*2048+ 411,   45*2048+ 412,   45*2048+ 413, 
  37*2048+ 414,    2*2048+ 415,    2*2048+ 416,   41*2048+ 417,   45*2048+ 418,   45*2048+ 419, 
   5*2048+ 420,    9*2048+ 421,   14*2048+ 422,   42*2048+ 423,   45*2048+ 424,   45*2048+ 425, 
  37*2048+ 426,   10*2048+ 427,    9*2048+ 428,    7*2048+ 429,   45*2048+ 430,   45*2048+ 431, 
  23*2048+ 432,    7*2048+ 433,   26*2048+ 434,   29*2048+ 435,   45*2048+ 436,   45*2048+ 437, 
  28*2048+ 438,   19*2048+ 439,    4*2048+ 440,    1*2048+ 441,   45*2048+ 442,   45*2048+ 443, 
  37*2048+ 444,   25*2048+ 445,   41*2048+ 446,   24*2048+ 447,   45*2048+ 448,   45*2048+ 449, 
  39*2048+ 450,   30*2048+ 451,    0*2048+ 452,   24*2048+ 453,   45*2048+ 454,   45*2048+ 455, 
  36*2048+ 456,   41*2048+ 457,   23*2048+ 458,   11*2048+ 459,   45*2048+ 460,   45*2048+ 461, 
   6*2048+ 462,   20*2048+ 463,   41*2048+ 464,   26*2048+ 465,   45*2048+ 466,   45*2048+ 467, 
  14*2048+ 468,    8*2048+ 469,   41*2048+ 470,    3*2048+ 471,   45*2048+ 472,   45*2048+ 473, 
   8*2048+ 474,    2*2048+ 475,   11*2048+ 476,    4*2048+ 477,   45*2048+ 478,   45*2048+ 479, 
  19*2048+ 480,   11*2048+ 481,   12*2048+ 482,    3*2048+ 483,   45*2048+ 484,   45*2048+ 485, 
   4*2048+ 486,    0*2048+ 487,   24*2048+ 488,   43*2048+ 489,   45*2048+ 490,   45*2048+ 491, 
  22*2048+ 492,   14*2048+ 493,   27*2048+ 494,   23*2048+ 495,   45*2048+ 496,   45*2048+ 497, 
  37*2048+ 498,   20*2048+ 499,    4*2048+ 500,   30*2048+ 501,   45*2048+ 502,   45*2048+ 503, 
  35*2048+ 504,   19*2048+ 505,   13*2048+ 506,   36*2048+ 507,   45*2048+ 508,   45*2048+ 509, 
   6*2048+ 510,   26*2048+ 511,   38*2048+ 512,   21*2048+ 513,   45*2048+ 514,   45*2048+ 515, 
  18*2048+ 516,   22*2048+ 517,   37*2048+ 518,    8*2048+ 519,   45*2048+ 520,   45*2048+ 521, 
  15*2048+ 522,    3*2048+ 523,   13*2048+ 524,    2*2048+ 525,   45*2048+ 526,   45*2048+ 527, 
  19*2048+ 528,    2*2048+ 529,   11*2048+ 530,   26*2048+ 531,   45*2048+ 532,   45*2048+ 533, 
  17*2048+ 534,   18*2048+ 535,   25*2048+ 536,    3*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
  42*2048+ 540,   15*2048+ 541,   33*2048+ 542,   14*2048+ 543,   45*2048+ 544,   45*2048+ 545, 
  39*2048+ 546,   13*2048+ 547,   43*2048+ 548,   21*2048+ 549,   45*2048+ 550,   45*2048+ 551, 
  44*2048+ 552,   36*2048+ 553,   37*2048+ 554,   24*2048+ 555,   45*2048+ 556,   45*2048+ 557, 
  26*2048+ 558,   37*2048+ 559,    4*2048+ 560,   18*2048+ 561,   45*2048+ 562,   45*2048+ 563, 
  35*2048+ 564,   35*2048+ 565,   33*2048+ 566,   27*2048+ 567,   45*2048+ 568,   45*2048+ 569, 
  43*2048+ 570,   33*2048+ 571,   42*2048+ 572,   36*2048+ 573,   45*2048+ 574,   45*2048+ 575, 
  37*2048+ 576,    2*2048+ 577,    2*2048+ 578,   41*2048+ 579,   45*2048+ 580,   45*2048+ 581, 
   5*2048+ 582,    9*2048+ 583,   14*2048+ 584,   42*2048+ 585,   45*2048+ 586,   45*2048+ 587, 
  37*2048+ 588,   10*2048+ 589,    9*2048+ 590,    7*2048+ 591,   45*2048+ 592,   45*2048+ 593, 
  23*2048+ 594,    7*2048+ 595,   26*2048+ 596,   29*2048+ 597,   45*2048+ 598,   45*2048+ 599, 
  28*2048+ 600,   19*2048+ 601,    4*2048+ 602,    1*2048+ 603,   45*2048+ 604,   45*2048+ 605, 
  37*2048+ 606,   25*2048+ 607,   41*2048+ 608,   24*2048+ 609,   45*2048+ 610,   45*2048+ 611, 
  25*2048+ 612,   39*2048+ 613,   30*2048+ 614,    0*2048+ 615,   45*2048+ 616,   45*2048+ 617, 
  36*2048+ 618,   41*2048+ 619,   23*2048+ 620,   11*2048+ 621,   45*2048+ 622,   45*2048+ 623, 
  27*2048+ 624,    6*2048+ 625,   20*2048+ 626,   41*2048+ 627,   45*2048+ 628,   45*2048+ 629, 
  14*2048+ 630,    8*2048+ 631,   41*2048+ 632,    3*2048+ 633,   45*2048+ 634,   45*2048+ 635, 
   8*2048+ 636,    2*2048+ 637,   11*2048+ 638,    4*2048+ 639,   45*2048+ 640,   45*2048+ 641, 
  13*2048+ 642,    4*2048+ 643,   19*2048+ 644,   11*2048+ 645,   45*2048+ 646,   45*2048+ 647, 
  25*2048+ 648,   44*2048+ 649,    4*2048+ 650,    0*2048+ 651,   45*2048+ 652,   45*2048+ 653, 
  28*2048+ 654,   24*2048+ 655,   22*2048+ 656,   14*2048+ 657,   45*2048+ 658,   45*2048+ 659, 
   5*2048+ 660,   31*2048+ 661,   37*2048+ 662,   20*2048+ 663,   45*2048+ 664,   45*2048+ 665, 
  35*2048+ 666,   19*2048+ 667,   13*2048+ 668,   36*2048+ 669,   45*2048+ 670,   45*2048+ 671, 
   6*2048+ 672,   26*2048+ 673,   38*2048+ 674,   21*2048+ 675,   45*2048+ 676,   45*2048+ 677, 
   9*2048+ 678,   18*2048+ 679,   22*2048+ 680,   37*2048+ 681,   45*2048+ 682,   45*2048+ 683, 
   4*2048+ 684,   14*2048+ 685,    3*2048+ 686,   15*2048+ 687,   45*2048+ 688,   45*2048+ 689, 
  19*2048+ 690,    2*2048+ 691,   11*2048+ 692,   26*2048+ 693,   45*2048+ 694,   45*2048+ 695, 
   4*2048+ 696,   17*2048+ 697,   18*2048+ 698,   25*2048+ 699,   45*2048+ 700,   45*2048+ 701, 
  15*2048+ 702,   42*2048+ 703,   15*2048+ 704,   33*2048+ 705,   45*2048+ 706,   45*2048+ 707, 
  39*2048+ 708,   13*2048+ 709,   43*2048+ 710,   21*2048+ 711,   45*2048+ 712,   45*2048+ 713, 
  25*2048+ 714,   44*2048+ 715,   36*2048+ 716,   37*2048+ 717,   45*2048+ 718,   45*2048+ 719, 
  26*2048+ 720,   37*2048+ 721,    4*2048+ 722,   18*2048+ 723,   45*2048+ 724,   45*2048+ 725, 
  35*2048+ 726,   35*2048+ 727,   33*2048+ 728,   27*2048+ 729,   45*2048+ 730,   45*2048+ 731, 
  43*2048+ 732,   33*2048+ 733,   42*2048+ 734,   36*2048+ 735,   45*2048+ 736,   45*2048+ 737, 
  42*2048+ 738,   37*2048+ 739,    2*2048+ 740,    2*2048+ 741,   45*2048+ 742,   45*2048+ 743, 
   5*2048+ 744,    9*2048+ 745,   14*2048+ 746,   42*2048+ 747,   45*2048+ 748,   45*2048+ 749, 
  37*2048+ 750,   10*2048+ 751,    9*2048+ 752,    7*2048+ 753,   45*2048+ 754,   45*2048+ 755, 
  30*2048+ 756,   23*2048+ 757,    7*2048+ 758,   26*2048+ 759,   45*2048+ 760,   45*2048+ 761, 
  28*2048+ 762,   19*2048+ 763,    4*2048+ 764,    1*2048+ 765,   45*2048+ 766,   45*2048+ 767, 
  37*2048+ 768,   25*2048+ 769,   41*2048+ 770,   24*2048+ 771,   45*2048+ 772,   45*2048+ 773, 
  25*2048+ 774,   39*2048+ 775,   30*2048+ 776,    0*2048+ 777,   45*2048+ 778,   45*2048+ 779, 
  12*2048+ 780,   36*2048+ 781,   41*2048+ 782,   23*2048+ 783,   45*2048+ 784,   45*2048+ 785, 
  27*2048+ 786,    6*2048+ 787,   20*2048+ 788,   41*2048+ 789,   45*2048+ 790,   45*2048+ 791, 
  14*2048+ 792,    8*2048+ 793,   41*2048+ 794,    3*2048+ 795,   45*2048+ 796,   45*2048+ 797, 
   8*2048+ 798,    2*2048+ 799,   11*2048+ 800,    4*2048+ 801,   45*2048+ 802,   45*2048+ 803, 
  13*2048+ 804,    4*2048+ 805,   19*2048+ 806,   11*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  25*2048+ 810,   44*2048+ 811,    4*2048+ 812,    0*2048+ 813,   45*2048+ 814,   45*2048+ 815, 
  28*2048+ 816,   24*2048+ 817,   22*2048+ 818,   14*2048+ 819,   45*2048+ 820,   45*2048+ 821, 
   5*2048+ 822,   31*2048+ 823,   37*2048+ 824,   20*2048+ 825,   45*2048+ 826,   45*2048+ 827, 
  37*2048+ 828,   35*2048+ 829,   19*2048+ 830,   13*2048+ 831,   45*2048+ 832,   45*2048+ 833, 
  39*2048+ 834,   22*2048+ 835,    6*2048+ 836,   26*2048+ 837,   45*2048+ 838,   45*2048+ 839, 
  38*2048+ 840,    9*2048+ 841,   18*2048+ 842,   22*2048+ 843,   45*2048+ 844,   45*2048+ 845, 
  16*2048+ 846,    4*2048+ 847,   14*2048+ 848,    3*2048+ 849,   45*2048+ 850,   45*2048+ 851, 
  27*2048+ 852,   19*2048+ 853,    2*2048+ 854,   11*2048+ 855,   45*2048+ 856,   45*2048+ 857, 
  26*2048+ 858,    4*2048+ 859,   17*2048+ 860,   18*2048+ 861,   45*2048+ 862,   45*2048+ 863, 
  34*2048+ 864,   15*2048+ 865,   42*2048+ 866,   15*2048+ 867,   45*2048+ 868,   45*2048+ 869, 
  39*2048+ 870,   13*2048+ 871,   43*2048+ 872,   21*2048+ 873,   45*2048+ 874,   45*2048+ 875, 
  25*2048+ 876,   44*2048+ 877,   36*2048+ 878,   37*2048+ 879,   45*2048+ 880,   45*2048+ 881, 
  26*2048+ 882,   37*2048+ 883,    4*2048+ 884,   18*2048+ 885,   45*2048+ 886,   45*2048+ 887, 
  35*2048+ 888,   35*2048+ 889,   33*2048+ 890,   27*2048+ 891,   45*2048+ 892,   45*2048+ 893, 
  43*2048+ 894,   33*2048+ 895,   42*2048+ 896,   36*2048+ 897,   45*2048+ 898,   45*2048+ 899, 
  42*2048+ 900,   37*2048+ 901,    2*2048+ 902,    2*2048+ 903,   45*2048+ 904,   45*2048+ 905, 
  43*2048+ 906,    5*2048+ 907,    9*2048+ 908,   14*2048+ 909,   45*2048+ 910,   45*2048+ 911, 
  37*2048+ 912,   10*2048+ 913,    9*2048+ 914,    7*2048+ 915,   45*2048+ 916,   45*2048+ 917, 
  27*2048+ 918,   30*2048+ 919,   23*2048+ 920,    7*2048+ 921,   45*2048+ 922,   45*2048+ 923, 
   2*2048+ 924,   28*2048+ 925,   19*2048+ 926,    4*2048+ 927,   45*2048+ 928,   45*2048+ 929, 
  37*2048+ 930,   25*2048+ 931,   41*2048+ 932,   24*2048+ 933,   45*2048+ 934,   45*2048+ 935, 
   1*2048+ 936,   25*2048+ 937,   39*2048+ 938,   30*2048+ 939,   45*2048+ 940,   45*2048+ 941, 
  12*2048+ 942,   36*2048+ 943,   41*2048+ 944,   23*2048+ 945,   45*2048+ 946,   45*2048+ 947, 
  42*2048+ 948,   27*2048+ 949,    6*2048+ 950,   20*2048+ 951,   45*2048+ 952,   45*2048+ 953, 
   4*2048+ 954,   14*2048+ 955,    8*2048+ 956,   41*2048+ 957,   45*2048+ 958,   45*2048+ 959, 
   8*2048+ 960,    2*2048+ 961,   11*2048+ 962,    4*2048+ 963,   45*2048+ 964,   45*2048+ 965, 
  13*2048+ 966,    4*2048+ 967,   19*2048+ 968,   11*2048+ 969,   45*2048+ 970,   45*2048+ 971, 
  25*2048+ 972,   44*2048+ 973,    4*2048+ 974,    0*2048+ 975,   45*2048+ 976,   45*2048+ 977, 
  28*2048+ 978,   24*2048+ 979,   22*2048+ 980,   14*2048+ 981,   45*2048+ 982,   45*2048+ 983, 
  21*2048+ 984,    5*2048+ 985,   31*2048+ 986,   37*2048+ 987,   45*2048+ 988,   45*2048+ 989, 
  37*2048+ 990,   35*2048+ 991,   19*2048+ 992,   13*2048+ 993,   45*2048+ 994,   45*2048+ 995, 
  39*2048+ 996,   22*2048+ 997,    6*2048+ 998,   26*2048+ 999,   45*2048+1000,   45*2048+1001, 
  38*2048+1002,    9*2048+1003,   18*2048+1004,   22*2048+1005,   45*2048+1006,   45*2048+1007, 
  16*2048+1008,    4*2048+1009,   14*2048+1010,    3*2048+1011,   45*2048+1012,   45*2048+1013, 
  27*2048+1014,   19*2048+1015,    2*2048+1016,   11*2048+1017,   45*2048+1018,   45*2048+1019, 
  26*2048+1020,    4*2048+1021,   17*2048+1022,   18*2048+1023,   45*2048+1024,   45*2048+1025, 
  34*2048+1026,   15*2048+1027,   42*2048+1028,   15*2048+1029,   45*2048+1030,   45*2048+1031, 
  22*2048+1032,   39*2048+1033,   13*2048+1034,   43*2048+1035,   45*2048+1036,   45*2048+1037, 
  38*2048+1038,   25*2048+1039,   44*2048+1040,   36*2048+1041,   45*2048+1042,   45*2048+1043, 
  19*2048+1044,   26*2048+1045,   37*2048+1046,    4*2048+1047,   45*2048+1048,   45*2048+1049, 
  28*2048+1050,   35*2048+1051,   35*2048+1052,   33*2048+1053,   45*2048+1054,   45*2048+1055, 
  43*2048+1056,   33*2048+1057,   42*2048+1058,   36*2048+1059,   45*2048+1060,   45*2048+1061, 
  42*2048+1062,   37*2048+1063,    2*2048+1064,    2*2048+1065,   45*2048+1066,   45*2048+1067, 
  15*2048+1068,   43*2048+1069,    5*2048+1070,    9*2048+1071,   45*2048+1072,   45*2048+1073, 
   8*2048+1074,   37*2048+1075,   10*2048+1076,    9*2048+1077,   45*2048+1078,   45*2048+1079, 
  27*2048+1080,   30*2048+1081,   23*2048+1082,    7*2048+1083,   45*2048+1084,   45*2048+1085, 
   5*2048+1086,    2*2048+1087,   28*2048+1088,   19*2048+1089,   45*2048+1090,   45*2048+1091, 
  25*2048+1092,   37*2048+1093,   25*2048+1094,   41*2048+1095,   45*2048+1096,   45*2048+1097, 
  31*2048+1098,    1*2048+1099,   25*2048+1100,   39*2048+1101,   45*2048+1102,   45*2048+1103, 
  12*2048+1104,   36*2048+1105,   41*2048+1106,   23*2048+1107,   45*2048+1108,   45*2048+1109, 
  42*2048+1110,   27*2048+1111,    6*2048+1112,   20*2048+1113,   45*2048+1114,   45*2048+1115, 
   4*2048+1116,   14*2048+1117,    8*2048+1118,   41*2048+1119,   45*2048+1120,   45*2048+1121, 
   5*2048+1122,    8*2048+1123,    2*2048+1124,   11*2048+1125,   45*2048+1126,   45*2048+1127, 
  13*2048+1128,    4*2048+1129,   19*2048+1130,   11*2048+1131,   45*2048+1132,   45*2048+1133, 
   1*2048+1134,   25*2048+1135,   44*2048+1136,    4*2048+1137,   45*2048+1138,   45*2048+1139, 
  28*2048+1140,   24*2048+1141,   22*2048+1142,   14*2048+1143,   45*2048+1144,   45*2048+1145, 
  21*2048+1146,    5*2048+1147,   31*2048+1148,   37*2048+1149,   45*2048+1150,   45*2048+1151, 
  37*2048+1152,   35*2048+1153,   19*2048+1154,   13*2048+1155,   45*2048+1156,   45*2048+1157, 
  39*2048+1158,   22*2048+1159,    6*2048+1160,   26*2048+1161,   45*2048+1162,   45*2048+1163, 
  23*2048+1164,   38*2048+1165,    9*2048+1166,   18*2048+1167,   45*2048+1168,   45*2048+1169, 
  16*2048+1170,    4*2048+1171,   14*2048+1172,    3*2048+1173,   45*2048+1174,   45*2048+1175, 
  27*2048+1176,   19*2048+1177,    2*2048+1178,   11*2048+1179,   45*2048+1180,   45*2048+1181, 
  26*2048+1182,    4*2048+1183,   17*2048+1184,   18*2048+1185,   45*2048+1186,   45*2048+1187, 
  34*2048+1188,   15*2048+1189,   42*2048+1190,   15*2048+1191,   45*2048+1192,   45*2048+1193, 
  44*2048+1194,   22*2048+1195,   39*2048+1196,   13*2048+1197,   45*2048+1198,   45*2048+1199, 
  37*2048+1200,   38*2048+1201,   25*2048+1202,   44*2048+1203,   45*2048+1204,   45*2048+1205, 
   5*2048+1206,   19*2048+1207,   26*2048+1208,   37*2048+1209,   45*2048+1210,   45*2048+1211, 
  28*2048+1212,   35*2048+1213,   35*2048+1214,   33*2048+1215,   45*2048+1216,   45*2048+1217, 
  43*2048+1218,   37*2048+1219,   43*2048+1220,   33*2048+1221,   45*2048+1222,   45*2048+1223, 
   3*2048+1224,   42*2048+1225,   37*2048+1226,    2*2048+1227,   45*2048+1228,   45*2048+1229, 
  15*2048+1230,   43*2048+1231,    5*2048+1232,    9*2048+1233,   45*2048+1234,   45*2048+1235, 
  10*2048+1236,    8*2048+1237,   37*2048+1238,   10*2048+1239,   45*2048+1240,   45*2048+1241, 
  27*2048+1242,   30*2048+1243,   23*2048+1244,    7*2048+1245,   45*2048+1246,   45*2048+1247, 
  20*2048+1248,    5*2048+1249,    2*2048+1250,   28*2048+1251,   45*2048+1252,   45*2048+1253, 
  42*2048+1254,   25*2048+1255,   37*2048+1256,   25*2048+1257,   45*2048+1258,   45*2048+1259, 
  31*2048+1260,    1*2048+1261,   25*2048+1262,   39*2048+1263,   45*2048+1264,   45*2048+1265, 
  12*2048+1266,   36*2048+1267,   41*2048+1268,   23*2048+1269,   45*2048+1270,   45*2048+1271, 
  21*2048+1272,   42*2048+1273,   27*2048+1274,    6*2048+1275,   45*2048+1276,   45*2048+1277, 
   4*2048+1278,   14*2048+1279,    8*2048+1280,   41*2048+1281,   45*2048+1282,   45*2048+1283, 
   3*2048+1284,   12*2048+1285,    5*2048+1286,    8*2048+1287,   45*2048+1288,   45*2048+1289, 
  13*2048+1290,    4*2048+1291,   19*2048+1292,   11*2048+1293,   45*2048+1294,   45*2048+1295, 

  45*2048+  24,   13*2048+  25,   45*2048+  26,   45*2048+  27, 
  45*2048+  33,   22*2048+  34,   45*2048+  35,   45*2048+  36, 
  39*2048+  87,   44*2048+  88,   45*2048+  89,   45*2048+  90, 
  11*2048+ 102,   43*2048+ 103,   45*2048+ 104,   45*2048+ 105, 
  45*2048+ 159,   13*2048+ 160,   45*2048+ 161,   45*2048+ 162, 
  45*2048+ 168,   22*2048+ 169,   45*2048+ 170,   45*2048+ 171, 
  39*2048+ 222,   44*2048+ 223,   45*2048+ 224,   45*2048+ 225, 
  11*2048+ 237,   43*2048+ 238,   45*2048+ 239,   45*2048+ 240, 
  45*2048+ 294,   13*2048+ 295,   45*2048+ 296,   45*2048+ 297, 
  45*2048+ 303,   22*2048+ 304,   45*2048+ 305,   45*2048+ 306, 
  45*2048+ 357,   39*2048+ 358,   45*2048+ 359,   45*2048+ 360, 
  44*2048+ 372,   11*2048+ 373,   45*2048+ 374,   45*2048+ 375, 
  45*2048+ 429,   13*2048+ 430,   45*2048+ 431,   45*2048+ 432, 
  45*2048+ 438,   22*2048+ 439,   45*2048+ 440,   45*2048+ 441, 
  40*2048+ 492,   45*2048+ 493,   45*2048+ 494,   45*2048+ 495, 
  12*2048+ 507,   44*2048+ 508,   45*2048+ 509,   45*2048+ 510, 
  45*2048+ 564,   13*2048+ 565,   45*2048+ 566,   45*2048+ 567, 
  45*2048+ 573,   22*2048+ 574,   45*2048+ 575,   45*2048+ 576, 
  40*2048+ 627,   45*2048+ 628,   45*2048+ 629,   45*2048+ 630, 
  12*2048+ 642,   44*2048+ 643,   45*2048+ 644,   45*2048+ 645, 
  45*2048+ 699,   13*2048+ 700,   45*2048+ 701,   45*2048+ 702, 
  45*2048+ 708,   22*2048+ 709,   45*2048+ 710,   45*2048+ 711, 
  40*2048+ 762,   45*2048+ 763,   45*2048+ 764,   45*2048+ 765, 
  12*2048+ 777,   44*2048+ 778,   45*2048+ 779,   45*2048+ 780, 
  14*2048+ 834,   45*2048+ 835,   45*2048+ 836,   45*2048+ 837, 
  45*2048+ 843,   22*2048+ 844,   45*2048+ 845,   45*2048+ 846, 
  40*2048+ 897,   45*2048+ 898,   45*2048+ 899,   45*2048+ 900, 
  12*2048+ 912,   44*2048+ 913,   45*2048+ 914,   45*2048+ 915, 
  14*2048+ 969,   45*2048+ 970,   45*2048+ 971,   45*2048+ 972, 
  45*2048+ 978,   22*2048+ 979,   45*2048+ 980,   45*2048+ 981, 
  40*2048+1032,   45*2048+1033,   45*2048+1034,   45*2048+1035, 
  12*2048+1047,   44*2048+1048,   45*2048+1049,   45*2048+1050, 
  45*2048+   0,   25*2048+   1,   27*2048+   2,   45*2048+   3,   44*2048+   4, 
  45*2048+  28,   29*2048+  29,   30*2048+  30,   45*2048+  31,   45*2048+  32, 
  45*2048+  37,   27*2048+  38,   39*2048+  39,   45*2048+  40,   45*2048+  41, 
  45*2048+  48,   10*2048+  49,   25*2048+  50,   45*2048+  51,   45*2048+  52, 
  45*2048+  53,   39*2048+  54,    0*2048+  55,   45*2048+  56,   45*2048+  57, 
  29*2048+  82,   19*2048+  83,   43*2048+  84,   45*2048+  85,   45*2048+  86, 
  32*2048+  97,   26*2048+  98,   10*2048+  99,   45*2048+ 100,   45*2048+ 101, 
  45*2048+ 112,   20*2048+ 113,   24*2048+ 114,   45*2048+ 115,   45*2048+ 116, 
  45*2048+ 123,   16*2048+ 124,   33*2048+ 125,   45*2048+ 126,   45*2048+ 127, 
  45*2048+ 135,   25*2048+ 136,   27*2048+ 137,   45*2048+ 138,   45*2048+ 139, 
  45*2048+ 163,   29*2048+ 164,   30*2048+ 165,   45*2048+ 166,   45*2048+ 167, 
  45*2048+ 172,   27*2048+ 173,   39*2048+ 174,   45*2048+ 175,   45*2048+ 176, 
  45*2048+ 183,   10*2048+ 184,   25*2048+ 185,   45*2048+ 186,   45*2048+ 187, 
  45*2048+ 188,   39*2048+ 189,    0*2048+ 190,   45*2048+ 191,   45*2048+ 192, 
  29*2048+ 217,   19*2048+ 218,   43*2048+ 219,   45*2048+ 220,   45*2048+ 221, 
  32*2048+ 232,   26*2048+ 233,   10*2048+ 234,   45*2048+ 235,   45*2048+ 236, 
  25*2048+ 247,   45*2048+ 248,   20*2048+ 249,   45*2048+ 250,   45*2048+ 251, 
  45*2048+ 258,   16*2048+ 259,   33*2048+ 260,   45*2048+ 261,   45*2048+ 262, 
  26*2048+ 270,   28*2048+ 271,   45*2048+ 272,   45*2048+ 273,   45*2048+ 274, 
  31*2048+ 298,   45*2048+ 299,   29*2048+ 300,   45*2048+ 301,   45*2048+ 302, 
  40*2048+ 307,   45*2048+ 308,   27*2048+ 309,   45*2048+ 310,   45*2048+ 311, 
  45*2048+ 318,   10*2048+ 319,   25*2048+ 320,   45*2048+ 321,   45*2048+ 322, 
  45*2048+ 323,   39*2048+ 324,    0*2048+ 325,   45*2048+ 326,   45*2048+ 327, 
  29*2048+ 352,   19*2048+ 353,   43*2048+ 354,   45*2048+ 355,   45*2048+ 356, 
  11*2048+ 367,   32*2048+ 368,   26*2048+ 369,   45*2048+ 370,   45*2048+ 371, 
  25*2048+ 382,   45*2048+ 383,   20*2048+ 384,   45*2048+ 385,   45*2048+ 386, 
  45*2048+ 393,   16*2048+ 394,   33*2048+ 395,   45*2048+ 396,   45*2048+ 397, 
  26*2048+ 405,   28*2048+ 406,   45*2048+ 407,   45*2048+ 408,   45*2048+ 409, 
  30*2048+ 433,   31*2048+ 434,   45*2048+ 435,   45*2048+ 436,   45*2048+ 437, 
  40*2048+ 442,   45*2048+ 443,   27*2048+ 444,   45*2048+ 445,   45*2048+ 446, 
  26*2048+ 453,   45*2048+ 454,   10*2048+ 455,   45*2048+ 456,   45*2048+ 457, 
  45*2048+ 458,   39*2048+ 459,    0*2048+ 460,   45*2048+ 461,   45*2048+ 462, 
  44*2048+ 487,   29*2048+ 488,   19*2048+ 489,   45*2048+ 490,   45*2048+ 491, 
  27*2048+ 502,   11*2048+ 503,   32*2048+ 504,   45*2048+ 505,   45*2048+ 506, 
  25*2048+ 517,   45*2048+ 518,   20*2048+ 519,   45*2048+ 520,   45*2048+ 521, 
  45*2048+ 528,   16*2048+ 529,   33*2048+ 530,   45*2048+ 531,   45*2048+ 532, 
  26*2048+ 540,   28*2048+ 541,   45*2048+ 542,   45*2048+ 543,   45*2048+ 544, 
  30*2048+ 568,   31*2048+ 569,   45*2048+ 570,   45*2048+ 571,   45*2048+ 572, 
  28*2048+ 577,   40*2048+ 578,   45*2048+ 579,   45*2048+ 580,   45*2048+ 581, 
  26*2048+ 588,   45*2048+ 589,   10*2048+ 590,   45*2048+ 591,   45*2048+ 592, 
  45*2048+ 593,   39*2048+ 594,    0*2048+ 595,   45*2048+ 596,   45*2048+ 597, 
  44*2048+ 622,   29*2048+ 623,   19*2048+ 624,   45*2048+ 625,   45*2048+ 626, 
  27*2048+ 637,   11*2048+ 638,   32*2048+ 639,   45*2048+ 640,   45*2048+ 641, 
  25*2048+ 652,   45*2048+ 653,   20*2048+ 654,   45*2048+ 655,   45*2048+ 656, 
  45*2048+ 663,   16*2048+ 664,   33*2048+ 665,   45*2048+ 666,   45*2048+ 667, 
  26*2048+ 675,   28*2048+ 676,   45*2048+ 677,   45*2048+ 678,   45*2048+ 679, 
  30*2048+ 703,   31*2048+ 704,   45*2048+ 705,   45*2048+ 706,   45*2048+ 707, 
  28*2048+ 712,   40*2048+ 713,   45*2048+ 714,   45*2048+ 715,   45*2048+ 716, 
  11*2048+ 723,   26*2048+ 724,   45*2048+ 725,   45*2048+ 726,   45*2048+ 727, 
   1*2048+ 728,   45*2048+ 729,   39*2048+ 730,   45*2048+ 731,   45*2048+ 732, 
  20*2048+ 757,   44*2048+ 758,   29*2048+ 759,   45*2048+ 760,   45*2048+ 761, 
  33*2048+ 772,   27*2048+ 773,   11*2048+ 774,   45*2048+ 775,   45*2048+ 776, 
  25*2048+ 787,   45*2048+ 788,   20*2048+ 789,   45*2048+ 790,   45*2048+ 791, 
  17*2048+ 798,   34*2048+ 799,   45*2048+ 800,   45*2048+ 801,   45*2048+ 802, 
  26*2048+ 810,   28*2048+ 811,   45*2048+ 812,   45*2048+ 813,   45*2048+ 814, 
  30*2048+ 838,   31*2048+ 839,   45*2048+ 840,   45*2048+ 841,   45*2048+ 842, 
  28*2048+ 847,   40*2048+ 848,   45*2048+ 849,   45*2048+ 850,   45*2048+ 851, 
  11*2048+ 858,   26*2048+ 859,   45*2048+ 860,   45*2048+ 861,   45*2048+ 862, 
   1*2048+ 863,   45*2048+ 864,   39*2048+ 865,   45*2048+ 866,   45*2048+ 867, 
  20*2048+ 892,   44*2048+ 893,   29*2048+ 894,   45*2048+ 895,   45*2048+ 896, 
  33*2048+ 907,   27*2048+ 908,   11*2048+ 909,   45*2048+ 910,   45*2048+ 911, 
  25*2048+ 922,   45*2048+ 923,   20*2048+ 924,   45*2048+ 925,   45*2048+ 926, 
  17*2048+ 933,   34*2048+ 934,   45*2048+ 935,   45*2048+ 936,   45*2048+ 937, 
  26*2048+ 945,   28*2048+ 946,   45*2048+ 947,   45*2048+ 948,   45*2048+ 949, 
  30*2048+ 973,   31*2048+ 974,   45*2048+ 975,   45*2048+ 976,   45*2048+ 977, 
  28*2048+ 982,   40*2048+ 983,   45*2048+ 984,   45*2048+ 985,   45*2048+ 986, 
  11*2048+ 993,   26*2048+ 994,   45*2048+ 995,   45*2048+ 996,   45*2048+ 997, 
  40*2048+ 998,    1*2048+ 999,   45*2048+1000,   45*2048+1001,   45*2048+1002, 
  30*2048+1027,   20*2048+1028,   44*2048+1029,   45*2048+1030,   45*2048+1031, 
  33*2048+1042,   27*2048+1043,   11*2048+1044,   45*2048+1045,   45*2048+1046, 
  21*2048+1057,   25*2048+1058,   45*2048+1059,   45*2048+1060,   45*2048+1061, 
  17*2048+1068,   34*2048+1069,   45*2048+1070,   45*2048+1071,   45*2048+1072, 
  45*2048+   5,   40*2048+   6,   16*2048+   7,   15*2048+   8,   45*2048+   9,   45*2048+  10, 
  35*2048+  18,   45*2048+  19,   13*2048+  20,   29*2048+  21,   45*2048+  22,   45*2048+  23, 
  45*2048+  42,   19*2048+  43,   39*2048+  44,   21*2048+  45,   45*2048+  46,   45*2048+  47, 
  45*2048+  58,    8*2048+  59,   33*2048+  60,   24*2048+  61,   45*2048+  62,   45*2048+  63, 
  44*2048+  64,   45*2048+  65,   41*2048+  66,   39*2048+  67,   45*2048+  68,   45*2048+  69, 
  45*2048+  70,   15*2048+  71,   38*2048+  72,   32*2048+  73,   45*2048+  74,   45*2048+  75, 
  45*2048+  76,   41*2048+  77,   29*2048+  78,   27*2048+  79,   45*2048+  80,   45*2048+  81, 
  21*2048+  91,   21*2048+  92,   37*2048+  93,   33*2048+  94,   45*2048+  95,   45*2048+  96, 
  45*2048+ 106,    6*2048+ 107,   22*2048+ 108,   19*2048+ 109,   45*2048+ 110,   45*2048+ 111, 
  21*2048+ 117,   45*2048+ 118,   23*2048+ 119,   12*2048+ 120,   45*2048+ 121,   45*2048+ 122, 
  45*2048+ 140,   40*2048+ 141,   16*2048+ 142,   15*2048+ 143,   45*2048+ 144,   45*2048+ 145, 
  30*2048+ 153,   35*2048+ 154,   45*2048+ 155,   13*2048+ 156,   45*2048+ 157,   45*2048+ 158, 
  22*2048+ 177,   45*2048+ 178,   19*2048+ 179,   39*2048+ 180,   45*2048+ 181,   45*2048+ 182, 
  45*2048+ 193,    8*2048+ 194,   33*2048+ 195,   24*2048+ 196,   45*2048+ 197,   45*2048+ 198, 
  44*2048+ 199,   45*2048+ 200,   41*2048+ 201,   39*2048+ 202,   45*2048+ 203,   45*2048+ 204, 
  33*2048+ 205,   45*2048+ 206,   15*2048+ 207,   38*2048+ 208,   45*2048+ 209,   45*2048+ 210, 
  28*2048+ 211,   45*2048+ 212,   41*2048+ 213,   29*2048+ 214,   45*2048+ 215,   45*2048+ 216, 
  34*2048+ 226,   21*2048+ 227,   21*2048+ 228,   37*2048+ 229,   45*2048+ 230,   45*2048+ 231, 
  20*2048+ 241,   45*2048+ 242,    6*2048+ 243,   22*2048+ 244,   45*2048+ 245,   45*2048+ 246, 
  21*2048+ 252,   45*2048+ 253,   23*2048+ 254,   12*2048+ 255,   45*2048+ 256,   45*2048+ 257, 
  45*2048+ 275,   40*2048+ 276,   16*2048+ 277,   15*2048+ 278,   45*2048+ 279,   45*2048+ 280, 
  30*2048+ 288,   35*2048+ 289,   45*2048+ 290,   13*2048+ 291,   45*2048+ 292,   45*2048+ 293, 
  22*2048+ 312,   45*2048+ 313,   19*2048+ 314,   39*2048+ 315,   45*2048+ 316,   45*2048+ 317, 
  25*2048+ 328,   45*2048+ 329,    8*2048+ 330,   33*2048+ 331,   45*2048+ 332,   45*2048+ 333, 
  40*2048+ 334,   44*2048+ 335,   45*2048+ 336,   41*2048+ 337,   45*2048+ 338,   45*2048+ 339, 
  39*2048+ 340,   33*2048+ 341,   45*2048+ 342,   15*2048+ 343,   45*2048+ 344,   45*2048+ 345, 
  28*2048+ 346,   45*2048+ 347,   41*2048+ 348,   29*2048+ 349,   45*2048+ 350,   45*2048+ 351, 
  22*2048+ 361,   38*2048+ 362,   34*2048+ 363,   21*2048+ 364,   45*2048+ 365,   45*2048+ 366, 
  20*2048+ 376,   45*2048+ 377,    6*2048+ 378,   22*2048+ 379,   45*2048+ 380,   45*2048+ 381, 
  21*2048+ 387,   45*2048+ 388,   23*2048+ 389,   12*2048+ 390,   45*2048+ 391,   45*2048+ 392, 
  16*2048+ 410,   45*2048+ 411,   40*2048+ 412,   16*2048+ 413,   45*2048+ 414,   45*2048+ 415, 
  30*2048+ 423,   35*2048+ 424,   45*2048+ 425,   13*2048+ 426,   45*2048+ 427,   45*2048+ 428, 
  22*2048+ 447,   45*2048+ 448,   19*2048+ 449,   39*2048+ 450,   45*2048+ 451,   45*2048+ 452, 
  25*2048+ 463,   45*2048+ 464,    8*2048+ 465,   33*2048+ 466,   45*2048+ 467,   45*2048+ 468, 
  40*2048+ 469,   44*2048+ 470,   45*2048+ 471,   41*2048+ 472,   45*2048+ 473,   45*2048+ 474, 
  39*2048+ 475,   33*2048+ 476,   45*2048+ 477,   15*2048+ 478,   45*2048+ 479,   45*2048+ 480, 
  30*2048+ 481,   28*2048+ 482,   45*2048+ 483,   41*2048+ 484,   45*2048+ 485,   45*2048+ 486, 
  22*2048+ 496,   38*2048+ 497,   34*2048+ 498,   21*2048+ 499,   45*2048+ 500,   45*2048+ 501, 
  20*2048+ 511,   45*2048+ 512,    6*2048+ 513,   22*2048+ 514,   45*2048+ 515,   45*2048+ 516, 
  13*2048+ 522,   21*2048+ 523,   45*2048+ 524,   23*2048+ 525,   45*2048+ 526,   45*2048+ 527, 
  17*2048+ 545,   16*2048+ 546,   45*2048+ 547,   40*2048+ 548,   45*2048+ 549,   45*2048+ 550, 
  30*2048+ 558,   35*2048+ 559,   45*2048+ 560,   13*2048+ 561,   45*2048+ 562,   45*2048+ 563, 
  22*2048+ 582,   45*2048+ 583,   19*2048+ 584,   39*2048+ 585,   45*2048+ 586,   45*2048+ 587, 
  25*2048+ 598,   45*2048+ 599,    8*2048+ 600,   33*2048+ 601,   45*2048+ 602,   45*2048+ 603, 
  42*2048+ 604,   40*2048+ 605,   44*2048+ 606,   45*2048+ 607,   45*2048+ 608,   45*2048+ 609, 
  39*2048+ 610,   33*2048+ 611,   45*2048+ 612,   15*2048+ 613,   45*2048+ 614,   45*2048+ 615, 
  30*2048+ 616,   28*2048+ 617,   45*2048+ 618,   41*2048+ 619,   45*2048+ 620,   45*2048+ 621, 
  22*2048+ 631,   38*2048+ 632,   34*2048+ 633,   21*2048+ 634,   45*2048+ 635,   45*2048+ 636, 
  23*2048+ 646,   20*2048+ 647,   45*2048+ 648,    6*2048+ 649,   45*2048+ 650,   45*2048+ 651, 
  13*2048+ 657,   21*2048+ 658,   45*2048+ 659,   23*2048+ 660,   45*2048+ 661,   45*2048+ 662, 
  41*2048+ 680,   17*2048+ 681,   16*2048+ 682,   45*2048+ 683,   45*2048+ 684,   45*2048+ 685, 
  14*2048+ 693,   30*2048+ 694,   35*2048+ 695,   45*2048+ 696,   45*2048+ 697,   45*2048+ 698, 
  22*2048+ 717,   45*2048+ 718,   19*2048+ 719,   39*2048+ 720,   45*2048+ 721,   45*2048+ 722, 
  25*2048+ 733,   45*2048+ 734,    8*2048+ 735,   33*2048+ 736,   45*2048+ 737,   45*2048+ 738, 
  42*2048+ 739,   40*2048+ 740,   44*2048+ 741,   45*2048+ 742,   45*2048+ 743,   45*2048+ 744, 
  39*2048+ 745,   33*2048+ 746,   45*2048+ 747,   15*2048+ 748,   45*2048+ 749,   45*2048+ 750, 
  30*2048+ 751,   28*2048+ 752,   45*2048+ 753,   41*2048+ 754,   45*2048+ 755,   45*2048+ 756, 
  22*2048+ 766,   22*2048+ 767,   38*2048+ 768,   34*2048+ 769,   45*2048+ 770,   45*2048+ 771, 
  23*2048+ 781,   20*2048+ 782,   45*2048+ 783,    6*2048+ 784,   45*2048+ 785,   45*2048+ 786, 
  13*2048+ 792,   21*2048+ 793,   45*2048+ 794,   23*2048+ 795,   45*2048+ 796,   45*2048+ 797, 
  41*2048+ 815,   17*2048+ 816,   16*2048+ 817,   45*2048+ 818,   45*2048+ 819,   45*2048+ 820, 
  14*2048+ 828,   30*2048+ 829,   35*2048+ 830,   45*2048+ 831,   45*2048+ 832,   45*2048+ 833, 
  20*2048+ 852,   40*2048+ 853,   22*2048+ 854,   45*2048+ 855,   45*2048+ 856,   45*2048+ 857, 
  25*2048+ 868,   45*2048+ 869,    8*2048+ 870,   33*2048+ 871,   45*2048+ 872,   45*2048+ 873, 
  42*2048+ 874,   40*2048+ 875,   44*2048+ 876,   45*2048+ 877,   45*2048+ 878,   45*2048+ 879, 
  39*2048+ 880,   33*2048+ 881,   45*2048+ 882,   15*2048+ 883,   45*2048+ 884,   45*2048+ 885, 
  42*2048+ 886,   30*2048+ 887,   28*2048+ 888,   45*2048+ 889,   45*2048+ 890,   45*2048+ 891, 
  22*2048+ 901,   22*2048+ 902,   38*2048+ 903,   34*2048+ 904,   45*2048+ 905,   45*2048+ 906, 
  23*2048+ 916,   20*2048+ 917,   45*2048+ 918,    6*2048+ 919,   45*2048+ 920,   45*2048+ 921, 
  13*2048+ 927,   21*2048+ 928,   45*2048+ 929,   23*2048+ 930,   45*2048+ 931,   45*2048+ 932, 
  41*2048+ 950,   17*2048+ 951,   16*2048+ 952,   45*2048+ 953,   45*2048+ 954,   45*2048+ 955, 
  14*2048+ 963,   30*2048+ 964,   35*2048+ 965,   45*2048+ 966,   45*2048+ 967,   45*2048+ 968, 
  20*2048+ 987,   40*2048+ 988,   22*2048+ 989,   45*2048+ 990,   45*2048+ 991,   45*2048+ 992, 
  34*2048+1003,   25*2048+1004,   45*2048+1005,    8*2048+1006,   45*2048+1007,   45*2048+1008, 
  42*2048+1009,   40*2048+1010,   44*2048+1011,   45*2048+1012,   45*2048+1013,   45*2048+1014, 
  16*2048+1015,   39*2048+1016,   33*2048+1017,   45*2048+1018,   45*2048+1019,   45*2048+1020, 
  42*2048+1021,   30*2048+1022,   28*2048+1023,   45*2048+1024,   45*2048+1025,   45*2048+1026, 
  22*2048+1036,   22*2048+1037,   38*2048+1038,   34*2048+1039,   45*2048+1040,   45*2048+1041, 
  23*2048+1051,   20*2048+1052,   45*2048+1053,    6*2048+1054,   45*2048+1055,   45*2048+1056, 
  13*2048+1062,   21*2048+1063,   45*2048+1064,   23*2048+1065,   45*2048+1066,   45*2048+1067, 
  31*2048+  11,   14*2048+  12,   45*2048+  13,   27*2048+  14,    5*2048+  15,   45*2048+  16,   45*2048+  17, 
  45*2048+ 128,   18*2048+ 129,   15*2048+ 130,   22*2048+ 131,   24*2048+ 132,   45*2048+ 133,   45*2048+ 134, 
  31*2048+ 146,   14*2048+ 147,   45*2048+ 148,   27*2048+ 149,    5*2048+ 150,   45*2048+ 151,   45*2048+ 152, 
  23*2048+ 263,   25*2048+ 264,   45*2048+ 265,   18*2048+ 266,   15*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
  31*2048+ 281,   14*2048+ 282,   45*2048+ 283,   27*2048+ 284,    5*2048+ 285,   45*2048+ 286,   45*2048+ 287, 
  23*2048+ 398,   25*2048+ 399,   45*2048+ 400,   18*2048+ 401,   15*2048+ 402,   45*2048+ 403,   45*2048+ 404, 
   6*2048+ 416,   31*2048+ 417,   14*2048+ 418,   45*2048+ 419,   27*2048+ 420,   45*2048+ 421,   45*2048+ 422, 
  23*2048+ 533,   25*2048+ 534,   45*2048+ 535,   18*2048+ 536,   15*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
   6*2048+ 551,   31*2048+ 552,   14*2048+ 553,   45*2048+ 554,   27*2048+ 555,   45*2048+ 556,   45*2048+ 557, 
  19*2048+ 668,   16*2048+ 669,   23*2048+ 670,   25*2048+ 671,   45*2048+ 672,   45*2048+ 673,   45*2048+ 674, 
   6*2048+ 686,   31*2048+ 687,   14*2048+ 688,   45*2048+ 689,   27*2048+ 690,   45*2048+ 691,   45*2048+ 692, 
  19*2048+ 803,   16*2048+ 804,   23*2048+ 805,   25*2048+ 806,   45*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
   6*2048+ 821,   31*2048+ 822,   14*2048+ 823,   45*2048+ 824,   27*2048+ 825,   45*2048+ 826,   45*2048+ 827, 
  19*2048+ 938,   16*2048+ 939,   23*2048+ 940,   25*2048+ 941,   45*2048+ 942,   45*2048+ 943,   45*2048+ 944, 
  28*2048+ 956,    6*2048+ 957,   31*2048+ 958,   14*2048+ 959,   45*2048+ 960,   45*2048+ 961,   45*2048+ 962, 
  19*2048+1073,   16*2048+1074,   23*2048+1075,   25*2048+1076,   45*2048+1077,   45*2048+1078,   45*2048+1079, 

  45*2048+   0,   30*2048+   1,   11*2048+   2,   15*2048+   3,   42*2048+   4,    0*2048+   5,   23*2048+   6,   18*2048+   7,   27*2048+   8,   45*2048+   9,   44*2048+  10, 
  30*2048+  11,   45*2048+  12,   16*2048+  13,    0*2048+  14,   31*2048+  15,   34*2048+  16,   10*2048+  17,    4*2048+  18,   16*2048+  19,   45*2048+  20,   45*2048+  21, 
  45*2048+  22,    1*2048+  23,   17*2048+  24,   42*2048+  25,   38*2048+  26,   13*2048+  27,   33*2048+  28,    5*2048+  29,   38*2048+  30,   45*2048+  31,   45*2048+  32, 
  40*2048+  33,    2*2048+  34,   45*2048+  35,    6*2048+  36,    4*2048+  37,   37*2048+  38,   23*2048+  39,   15*2048+  40,   34*2048+  41,   45*2048+  42,   45*2048+  43, 
  45*2048+  44,   12*2048+  45,   41*2048+  46,   36*2048+  47,   25*2048+  48,    5*2048+  49,   21*2048+  50,   32*2048+  51,   29*2048+  52,   45*2048+  53,   45*2048+  54, 
  12*2048+  55,   45*2048+  56,   33*2048+  57,   41*2048+  58,   37*2048+  59,   11*2048+  60,   44*2048+  61,   26*2048+  62,   24*2048+  63,   45*2048+  64,   45*2048+  65, 
  45*2048+  66,    8*2048+  67,   35*2048+  68,   26*2048+  69,   35*2048+  70,   14*2048+  71,   18*2048+  72,   29*2048+  73,    8*2048+  74,   45*2048+  75,   45*2048+  76, 
  29*2048+  77,   45*2048+  78,   23*2048+  79,    5*2048+  80,   39*2048+  81,   22*2048+  82,   26*2048+  83,   10*2048+  84,   15*2048+  85,   45*2048+  86,   45*2048+  87, 
  45*2048+  88,   15*2048+  89,   11*2048+  90,   20*2048+  91,   15*2048+  92,   18*2048+  93,    6*2048+  94,   24*2048+  95,    5*2048+  96,   45*2048+  97,   45*2048+  98, 
  45*2048+  99,   16*2048+ 100,   24*2048+ 101,   22*2048+ 102,    9*2048+ 103,   12*2048+ 104,    7*2048+ 105,    3*2048+ 106,   18*2048+ 107,   45*2048+ 108,   45*2048+ 109, 
  14*2048+ 110,   45*2048+ 111,   19*2048+ 112,    3*2048+ 113,   27*2048+ 114,   21*2048+ 115,   21*2048+ 116,   31*2048+ 117,    1*2048+ 118,   45*2048+ 119,   45*2048+ 120, 
  39*2048+ 121,   45*2048+ 122,   12*2048+ 123,   28*2048+ 124,   33*2048+ 125,   17*2048+ 126,   30*2048+ 127,   25*2048+ 128,   28*2048+ 129,   45*2048+ 130,   45*2048+ 131, 
  45*2048+ 132,   11*2048+ 133,   32*2048+ 134,   35*2048+ 135,   43*2048+ 136,   29*2048+ 137,   24*2048+ 138,    5*2048+ 139,    0*2048+ 140,   45*2048+ 141,   45*2048+ 142, 
  45*2048+ 143,   20*2048+ 144,   43*2048+ 145,   33*2048+ 146,   43*2048+ 147,    4*2048+ 148,   37*2048+ 149,   17*2048+ 150,   17*2048+ 151,   45*2048+ 152,   45*2048+ 153, 
   3*2048+ 154,   45*2048+ 155,   20*2048+ 156,   42*2048+ 157,   12*2048+ 158,   43*2048+ 159,   25*2048+ 160,   17*2048+ 161,   15*2048+ 162,   45*2048+ 163,   45*2048+ 164, 
  45*2048+ 165,    3*2048+ 166,    5*2048+ 167,   36*2048+ 168,   21*2048+ 169,   20*2048+ 170,    7*2048+ 171,    9*2048+ 172,   39*2048+ 173,   45*2048+ 174,   45*2048+ 175, 
  40*2048+ 176,   45*2048+ 177,    1*2048+ 178,   28*2048+ 179,   12*2048+ 180,    3*2048+ 181,   15*2048+ 182,   13*2048+ 183,   17*2048+ 184,   45*2048+ 185,   45*2048+ 186, 
   5*2048+ 187,   11*2048+ 188,   45*2048+ 189,   43*2048+ 190,   36*2048+ 191,   19*2048+ 192,    3*2048+ 193,   24*2048+ 194,   36*2048+ 195,   45*2048+ 196,   45*2048+ 197, 
  45*2048+ 198,   30*2048+ 199,   11*2048+ 200,   15*2048+ 201,   42*2048+ 202,    0*2048+ 203,   23*2048+ 204,   18*2048+ 205,   27*2048+ 206,   45*2048+ 207,   45*2048+ 208, 
  30*2048+ 209,   45*2048+ 210,   16*2048+ 211,    0*2048+ 212,   31*2048+ 213,   34*2048+ 214,   10*2048+ 215,    4*2048+ 216,   16*2048+ 217,   45*2048+ 218,   45*2048+ 219, 
  39*2048+ 220,   45*2048+ 221,    1*2048+ 222,   17*2048+ 223,   42*2048+ 224,   38*2048+ 225,   13*2048+ 226,   33*2048+ 227,    5*2048+ 228,   45*2048+ 229,   45*2048+ 230, 
  35*2048+ 231,   40*2048+ 232,    2*2048+ 233,   45*2048+ 234,    6*2048+ 235,    4*2048+ 236,   37*2048+ 237,   23*2048+ 238,   15*2048+ 239,   45*2048+ 240,   45*2048+ 241, 
  30*2048+ 242,   45*2048+ 243,   12*2048+ 244,   41*2048+ 245,   36*2048+ 246,   25*2048+ 247,    5*2048+ 248,   21*2048+ 249,   32*2048+ 250,   45*2048+ 251,   45*2048+ 252, 
  27*2048+ 253,   25*2048+ 254,   12*2048+ 255,   45*2048+ 256,   33*2048+ 257,   41*2048+ 258,   37*2048+ 259,   11*2048+ 260,   44*2048+ 261,   45*2048+ 262,   45*2048+ 263, 
  30*2048+ 264,    9*2048+ 265,   45*2048+ 266,    8*2048+ 267,   35*2048+ 268,   26*2048+ 269,   35*2048+ 270,   14*2048+ 271,   18*2048+ 272,   45*2048+ 273,   45*2048+ 274, 
  16*2048+ 275,   29*2048+ 276,   45*2048+ 277,   23*2048+ 278,    5*2048+ 279,   39*2048+ 280,   22*2048+ 281,   26*2048+ 282,   10*2048+ 283,   45*2048+ 284,   45*2048+ 285, 
  25*2048+ 286,    6*2048+ 287,   45*2048+ 288,   15*2048+ 289,   11*2048+ 290,   20*2048+ 291,   15*2048+ 292,   18*2048+ 293,    6*2048+ 294,   45*2048+ 295,   45*2048+ 296, 
  45*2048+ 297,   16*2048+ 298,   24*2048+ 299,   22*2048+ 300,    9*2048+ 301,   12*2048+ 302,    7*2048+ 303,    3*2048+ 304,   18*2048+ 305,   45*2048+ 306,   45*2048+ 307, 
  14*2048+ 308,   45*2048+ 309,   19*2048+ 310,    3*2048+ 311,   27*2048+ 312,   21*2048+ 313,   21*2048+ 314,   31*2048+ 315,    1*2048+ 316,   45*2048+ 317,   45*2048+ 318, 
  26*2048+ 319,   29*2048+ 320,   39*2048+ 321,   45*2048+ 322,   12*2048+ 323,   28*2048+ 324,   33*2048+ 325,   17*2048+ 326,   30*2048+ 327,   45*2048+ 328,   45*2048+ 329, 
  45*2048+ 330,   11*2048+ 331,   32*2048+ 332,   35*2048+ 333,   43*2048+ 334,   29*2048+ 335,   24*2048+ 336,    5*2048+ 337,    0*2048+ 338,   45*2048+ 339,   45*2048+ 340, 
  18*2048+ 341,   45*2048+ 342,   20*2048+ 343,   43*2048+ 344,   33*2048+ 345,   43*2048+ 346,    4*2048+ 347,   37*2048+ 348,   17*2048+ 349,   45*2048+ 350,   45*2048+ 351, 
   3*2048+ 352,   45*2048+ 353,   20*2048+ 354,   42*2048+ 355,   12*2048+ 356,   43*2048+ 357,   25*2048+ 358,   17*2048+ 359,   15*2048+ 360,   45*2048+ 361,   45*2048+ 362, 
  45*2048+ 363,    3*2048+ 364,    5*2048+ 365,   36*2048+ 366,   21*2048+ 367,   20*2048+ 368,    7*2048+ 369,    9*2048+ 370,   39*2048+ 371,   45*2048+ 372,   45*2048+ 373, 
  40*2048+ 374,   45*2048+ 375,    1*2048+ 376,   28*2048+ 377,   12*2048+ 378,    3*2048+ 379,   15*2048+ 380,   13*2048+ 381,   17*2048+ 382,   45*2048+ 383,   45*2048+ 384, 
   5*2048+ 385,   11*2048+ 386,   45*2048+ 387,   43*2048+ 388,   36*2048+ 389,   19*2048+ 390,    3*2048+ 391,   24*2048+ 392,   36*2048+ 393,   45*2048+ 394,   45*2048+ 395, 
  45*2048+ 396,   30*2048+ 397,   11*2048+ 398,   15*2048+ 399,   42*2048+ 400,    0*2048+ 401,   23*2048+ 402,   18*2048+ 403,   27*2048+ 404,   45*2048+ 405,   45*2048+ 406, 
   5*2048+ 407,   17*2048+ 408,   30*2048+ 409,   45*2048+ 410,   16*2048+ 411,    0*2048+ 412,   31*2048+ 413,   34*2048+ 414,   10*2048+ 415,   45*2048+ 416,   45*2048+ 417, 
  34*2048+ 418,    6*2048+ 419,   39*2048+ 420,   45*2048+ 421,    1*2048+ 422,   17*2048+ 423,   42*2048+ 424,   38*2048+ 425,   13*2048+ 426,   45*2048+ 427,   45*2048+ 428, 
  16*2048+ 429,   35*2048+ 430,   40*2048+ 431,    2*2048+ 432,   45*2048+ 433,    6*2048+ 434,    4*2048+ 435,   37*2048+ 436,   23*2048+ 437,   45*2048+ 438,   45*2048+ 439, 
  30*2048+ 440,   45*2048+ 441,   12*2048+ 442,   41*2048+ 443,   36*2048+ 444,   25*2048+ 445,    5*2048+ 446,   21*2048+ 447,   32*2048+ 448,   45*2048+ 449,   45*2048+ 450, 
  27*2048+ 451,   25*2048+ 452,   12*2048+ 453,   45*2048+ 454,   33*2048+ 455,   41*2048+ 456,   37*2048+ 457,   11*2048+ 458,   44*2048+ 459,   45*2048+ 460,   45*2048+ 461, 
  15*2048+ 462,   19*2048+ 463,   30*2048+ 464,    9*2048+ 465,   45*2048+ 466,    8*2048+ 467,   35*2048+ 468,   26*2048+ 469,   35*2048+ 470,   45*2048+ 471,   45*2048+ 472, 
  11*2048+ 473,   16*2048+ 474,   29*2048+ 475,   45*2048+ 476,   23*2048+ 477,    5*2048+ 478,   39*2048+ 479,   22*2048+ 480,   26*2048+ 481,   45*2048+ 482,   45*2048+ 483, 
   7*2048+ 484,   25*2048+ 485,    6*2048+ 486,   45*2048+ 487,   15*2048+ 488,   11*2048+ 489,   20*2048+ 490,   15*2048+ 491,   18*2048+ 492,   45*2048+ 493,   45*2048+ 494, 
  45*2048+ 495,   16*2048+ 496,   24*2048+ 497,   22*2048+ 498,    9*2048+ 499,   12*2048+ 500,    7*2048+ 501,    3*2048+ 502,   18*2048+ 503,   45*2048+ 504,   45*2048+ 505, 
   2*2048+ 506,   14*2048+ 507,   45*2048+ 508,   19*2048+ 509,    3*2048+ 510,   27*2048+ 511,   21*2048+ 512,   21*2048+ 513,   31*2048+ 514,   45*2048+ 515,   45*2048+ 516, 
  31*2048+ 517,   26*2048+ 518,   29*2048+ 519,   39*2048+ 520,   45*2048+ 521,   12*2048+ 522,   28*2048+ 523,   33*2048+ 524,   17*2048+ 525,   45*2048+ 526,   45*2048+ 527, 
  30*2048+ 528,   25*2048+ 529,    6*2048+ 530,    1*2048+ 531,   45*2048+ 532,   11*2048+ 533,   32*2048+ 534,   35*2048+ 535,   43*2048+ 536,   45*2048+ 537,   45*2048+ 538, 
   5*2048+ 539,   38*2048+ 540,   18*2048+ 541,   18*2048+ 542,   45*2048+ 543,   20*2048+ 544,   43*2048+ 545,   33*2048+ 546,   43*2048+ 547,   45*2048+ 548,   45*2048+ 549, 
   3*2048+ 550,   45*2048+ 551,   20*2048+ 552,   42*2048+ 553,   12*2048+ 554,   43*2048+ 555,   25*2048+ 556,   17*2048+ 557,   15*2048+ 558,   45*2048+ 559,   45*2048+ 560, 
  40*2048+ 561,   45*2048+ 562,    3*2048+ 563,    5*2048+ 564,   36*2048+ 565,   21*2048+ 566,   20*2048+ 567,    7*2048+ 568,    9*2048+ 569,   45*2048+ 570,   45*2048+ 571, 
  18*2048+ 572,   40*2048+ 573,   45*2048+ 574,    1*2048+ 575,   28*2048+ 576,   12*2048+ 577,    3*2048+ 578,   15*2048+ 579,   13*2048+ 580,   45*2048+ 581,   45*2048+ 582, 
  37*2048+ 583,    5*2048+ 584,   11*2048+ 585,   45*2048+ 586,   43*2048+ 587,   36*2048+ 588,   19*2048+ 589,    3*2048+ 590,   24*2048+ 591,   45*2048+ 592,   45*2048+ 593, 
  28*2048+ 594,   45*2048+ 595,   30*2048+ 596,   11*2048+ 597,   15*2048+ 598,   42*2048+ 599,    0*2048+ 600,   23*2048+ 601,   18*2048+ 602,   45*2048+ 603,   45*2048+ 604, 
  11*2048+ 605,    5*2048+ 606,   17*2048+ 607,   30*2048+ 608,   45*2048+ 609,   16*2048+ 610,    0*2048+ 611,   31*2048+ 612,   34*2048+ 613,   45*2048+ 614,   45*2048+ 615, 
  34*2048+ 616,    6*2048+ 617,   39*2048+ 618,   45*2048+ 619,    1*2048+ 620,   17*2048+ 621,   42*2048+ 622,   38*2048+ 623,   13*2048+ 624,   45*2048+ 625,   45*2048+ 626, 
  24*2048+ 627,   16*2048+ 628,   35*2048+ 629,   40*2048+ 630,    2*2048+ 631,   45*2048+ 632,    6*2048+ 633,    4*2048+ 634,   37*2048+ 635,   45*2048+ 636,   45*2048+ 637, 
  33*2048+ 638,   30*2048+ 639,   45*2048+ 640,   12*2048+ 641,   41*2048+ 642,   36*2048+ 643,   25*2048+ 644,    5*2048+ 645,   21*2048+ 646,   45*2048+ 647,   45*2048+ 648, 
  12*2048+ 649,   45*2048+ 650,   27*2048+ 651,   25*2048+ 652,   12*2048+ 653,   45*2048+ 654,   33*2048+ 655,   41*2048+ 656,   37*2048+ 657,   45*2048+ 658,   45*2048+ 659, 
  36*2048+ 660,   15*2048+ 661,   19*2048+ 662,   30*2048+ 663,    9*2048+ 664,   45*2048+ 665,    8*2048+ 666,   35*2048+ 667,   26*2048+ 668,   45*2048+ 669,   45*2048+ 670, 
  27*2048+ 671,   11*2048+ 672,   16*2048+ 673,   29*2048+ 674,   45*2048+ 675,   23*2048+ 676,    5*2048+ 677,   39*2048+ 678,   22*2048+ 679,   45*2048+ 680,   45*2048+ 681, 
  19*2048+ 682,    7*2048+ 683,   25*2048+ 684,    6*2048+ 685,   45*2048+ 686,   15*2048+ 687,   11*2048+ 688,   20*2048+ 689,   15*2048+ 690,   45*2048+ 691,   45*2048+ 692, 
  19*2048+ 693,   45*2048+ 694,   16*2048+ 695,   24*2048+ 696,   22*2048+ 697,    9*2048+ 698,   12*2048+ 699,    7*2048+ 700,    3*2048+ 701,   45*2048+ 702,   45*2048+ 703, 
  32*2048+ 704,    2*2048+ 705,   14*2048+ 706,   45*2048+ 707,   19*2048+ 708,    3*2048+ 709,   27*2048+ 710,   21*2048+ 711,   21*2048+ 712,   45*2048+ 713,   45*2048+ 714, 
  31*2048+ 715,   26*2048+ 716,   29*2048+ 717,   39*2048+ 718,   45*2048+ 719,   12*2048+ 720,   28*2048+ 721,   33*2048+ 722,   17*2048+ 723,   45*2048+ 724,   45*2048+ 725, 
  44*2048+ 726,   30*2048+ 727,   25*2048+ 728,    6*2048+ 729,    1*2048+ 730,   45*2048+ 731,   11*2048+ 732,   32*2048+ 733,   35*2048+ 734,   45*2048+ 735,   45*2048+ 736, 
  44*2048+ 737,    5*2048+ 738,   38*2048+ 739,   18*2048+ 740,   18*2048+ 741,   45*2048+ 742,   20*2048+ 743,   43*2048+ 744,   33*2048+ 745,   45*2048+ 746,   45*2048+ 747, 
  18*2048+ 748,   16*2048+ 749,    3*2048+ 750,   45*2048+ 751,   20*2048+ 752,   42*2048+ 753,   12*2048+ 754,   43*2048+ 755,   25*2048+ 756,   45*2048+ 757,   45*2048+ 758, 
  10*2048+ 759,   40*2048+ 760,   45*2048+ 761,    3*2048+ 762,    5*2048+ 763,   36*2048+ 764,   21*2048+ 765,   20*2048+ 766,    7*2048+ 767,   45*2048+ 768,   45*2048+ 769, 
  14*2048+ 770,   18*2048+ 771,   40*2048+ 772,   45*2048+ 773,    1*2048+ 774,   28*2048+ 775,   12*2048+ 776,    3*2048+ 777,   15*2048+ 778,   45*2048+ 779,   45*2048+ 780, 
  25*2048+ 781,   37*2048+ 782,    5*2048+ 783,   11*2048+ 784,   45*2048+ 785,   43*2048+ 786,   36*2048+ 787,   19*2048+ 788,    3*2048+ 789,   45*2048+ 790,   45*2048+ 791, 
  24*2048+ 792,   19*2048+ 793,   28*2048+ 794,   45*2048+ 795,   30*2048+ 796,   11*2048+ 797,   15*2048+ 798,   42*2048+ 799,    0*2048+ 800,   45*2048+ 801,   45*2048+ 802, 
  35*2048+ 803,   11*2048+ 804,    5*2048+ 805,   17*2048+ 806,   30*2048+ 807,   45*2048+ 808,   16*2048+ 809,    0*2048+ 810,   31*2048+ 811,   45*2048+ 812,   45*2048+ 813, 
  34*2048+ 814,    6*2048+ 815,   39*2048+ 816,   45*2048+ 817,    1*2048+ 818,   17*2048+ 819,   42*2048+ 820,   38*2048+ 821,   13*2048+ 822,   45*2048+ 823,   45*2048+ 824, 
  24*2048+ 825,   16*2048+ 826,   35*2048+ 827,   40*2048+ 828,    2*2048+ 829,   45*2048+ 830,    6*2048+ 831,    4*2048+ 832,   37*2048+ 833,   45*2048+ 834,   45*2048+ 835, 
   6*2048+ 836,   22*2048+ 837,   33*2048+ 838,   30*2048+ 839,   45*2048+ 840,   12*2048+ 841,   41*2048+ 842,   36*2048+ 843,   25*2048+ 844,   45*2048+ 845,   45*2048+ 846, 
  12*2048+ 847,   45*2048+ 848,   27*2048+ 849,   25*2048+ 850,   12*2048+ 851,   45*2048+ 852,   33*2048+ 853,   41*2048+ 854,   37*2048+ 855,   45*2048+ 856,   45*2048+ 857, 
  36*2048+ 858,   27*2048+ 859,   36*2048+ 860,   15*2048+ 861,   19*2048+ 862,   30*2048+ 863,    9*2048+ 864,   45*2048+ 865,    8*2048+ 866,   45*2048+ 867,   45*2048+ 868, 
  23*2048+ 869,   27*2048+ 870,   11*2048+ 871,   16*2048+ 872,   29*2048+ 873,   45*2048+ 874,   23*2048+ 875,    5*2048+ 876,   39*2048+ 877,   45*2048+ 878,   45*2048+ 879, 
  19*2048+ 880,    7*2048+ 881,   25*2048+ 882,    6*2048+ 883,   45*2048+ 884,   15*2048+ 885,   11*2048+ 886,   20*2048+ 887,   15*2048+ 888,   45*2048+ 889,   45*2048+ 890, 
   8*2048+ 891,    4*2048+ 892,   19*2048+ 893,   45*2048+ 894,   16*2048+ 895,   24*2048+ 896,   22*2048+ 897,    9*2048+ 898,   12*2048+ 899,   45*2048+ 900,   45*2048+ 901, 
  22*2048+ 902,   32*2048+ 903,    2*2048+ 904,   14*2048+ 905,   45*2048+ 906,   19*2048+ 907,    3*2048+ 908,   27*2048+ 909,   21*2048+ 910,   45*2048+ 911,   45*2048+ 912, 
  18*2048+ 913,   31*2048+ 914,   26*2048+ 915,   29*2048+ 916,   39*2048+ 917,   45*2048+ 918,   12*2048+ 919,   28*2048+ 920,   33*2048+ 921,   45*2048+ 922,   45*2048+ 923, 
  36*2048+ 924,   44*2048+ 925,   30*2048+ 926,   25*2048+ 927,    6*2048+ 928,    1*2048+ 929,   45*2048+ 930,   11*2048+ 931,   32*2048+ 932,   45*2048+ 933,   45*2048+ 934, 
  44*2048+ 935,    5*2048+ 936,   38*2048+ 937,   18*2048+ 938,   18*2048+ 939,   45*2048+ 940,   20*2048+ 941,   43*2048+ 942,   33*2048+ 943,   45*2048+ 944,   45*2048+ 945, 
  18*2048+ 946,   16*2048+ 947,    3*2048+ 948,   45*2048+ 949,   20*2048+ 950,   42*2048+ 951,   12*2048+ 952,   43*2048+ 953,   25*2048+ 954,   45*2048+ 955,   45*2048+ 956, 
  21*2048+ 957,    8*2048+ 958,   10*2048+ 959,   40*2048+ 960,   45*2048+ 961,    3*2048+ 962,    5*2048+ 963,   36*2048+ 964,   21*2048+ 965,   45*2048+ 966,   45*2048+ 967, 
  14*2048+ 968,   18*2048+ 969,   40*2048+ 970,   45*2048+ 971,    1*2048+ 972,   28*2048+ 973,   12*2048+ 974,    3*2048+ 975,   15*2048+ 976,   45*2048+ 977,   45*2048+ 978, 
   4*2048+ 979,   25*2048+ 980,   37*2048+ 981,    5*2048+ 982,   11*2048+ 983,   45*2048+ 984,   43*2048+ 985,   36*2048+ 986,   19*2048+ 987,   45*2048+ 988,   45*2048+ 989, 
   1*2048+ 990,   24*2048+ 991,   19*2048+ 992,   28*2048+ 993,   45*2048+ 994,   30*2048+ 995,   11*2048+ 996,   15*2048+ 997,   42*2048+ 998,   45*2048+ 999,   45*2048+1000, 
  35*2048+1001,   11*2048+1002,    5*2048+1003,   17*2048+1004,   30*2048+1005,   45*2048+1006,   16*2048+1007,    0*2048+1008,   31*2048+1009,   45*2048+1010,   45*2048+1011, 
  39*2048+1012,   14*2048+1013,   34*2048+1014,    6*2048+1015,   39*2048+1016,   45*2048+1017,    1*2048+1018,   17*2048+1019,   42*2048+1020,   45*2048+1021,   45*2048+1022, 
  24*2048+1023,   16*2048+1024,   35*2048+1025,   40*2048+1026,    2*2048+1027,   45*2048+1028,    6*2048+1029,    4*2048+1030,   37*2048+1031,   45*2048+1032,   45*2048+1033, 
  37*2048+1034,   26*2048+1035,    6*2048+1036,   22*2048+1037,   33*2048+1038,   30*2048+1039,   45*2048+1040,   12*2048+1041,   41*2048+1042,   45*2048+1043,   45*2048+1044, 
  12*2048+1045,   45*2048+1046,   27*2048+1047,   25*2048+1048,   12*2048+1049,   45*2048+1050,   33*2048+1051,   41*2048+1052,   37*2048+1053,   45*2048+1054,   45*2048+1055, 
  36*2048+1056,   27*2048+1057,   36*2048+1058,   15*2048+1059,   19*2048+1060,   30*2048+1061,    9*2048+1062,   45*2048+1063,    8*2048+1064,   45*2048+1065,   45*2048+1066, 
   6*2048+1067,   40*2048+1068,   23*2048+1069,   27*2048+1070,   11*2048+1071,   16*2048+1072,   29*2048+1073,   45*2048+1074,   23*2048+1075,   45*2048+1076,   45*2048+1077, 
  19*2048+1078,    7*2048+1079,   25*2048+1080,    6*2048+1081,   45*2048+1082,   15*2048+1083,   11*2048+1084,   20*2048+1085,   15*2048+1086,   45*2048+1087,   45*2048+1088, 
  10*2048+1089,   13*2048+1090,    8*2048+1091,    4*2048+1092,   19*2048+1093,   45*2048+1094,   16*2048+1095,   24*2048+1096,   22*2048+1097,   45*2048+1098,   45*2048+1099, 
  22*2048+1100,   22*2048+1101,   32*2048+1102,    2*2048+1103,   14*2048+1104,   45*2048+1105,   19*2048+1106,    3*2048+1107,   27*2048+1108,   45*2048+1109,   45*2048+1110, 
  18*2048+1111,   31*2048+1112,   26*2048+1113,   29*2048+1114,   39*2048+1115,   45*2048+1116,   12*2048+1117,   28*2048+1118,   33*2048+1119,   45*2048+1120,   45*2048+1121, 
  36*2048+1122,   44*2048+1123,   30*2048+1124,   25*2048+1125,    6*2048+1126,    1*2048+1127,   45*2048+1128,   11*2048+1129,   32*2048+1130,   45*2048+1131,   45*2048+1132, 
  44*2048+1133,    5*2048+1134,   38*2048+1135,   18*2048+1136,   18*2048+1137,   45*2048+1138,   20*2048+1139,   43*2048+1140,   33*2048+1141,   45*2048+1142,   45*2048+1143, 
  26*2048+1144,   18*2048+1145,   16*2048+1146,    3*2048+1147,   45*2048+1148,   20*2048+1149,   42*2048+1150,   12*2048+1151,   43*2048+1152,   45*2048+1153,   45*2048+1154, 
  37*2048+1155,   22*2048+1156,   21*2048+1157,    8*2048+1158,   10*2048+1159,   40*2048+1160,   45*2048+1161,    3*2048+1162,    5*2048+1163,   45*2048+1164,   45*2048+1165, 
  16*2048+1166,   14*2048+1167,   18*2048+1168,   40*2048+1169,   45*2048+1170,    1*2048+1171,   28*2048+1172,   12*2048+1173,    3*2048+1174,   45*2048+1175,   45*2048+1176, 
  20*2048+1177,    4*2048+1178,   25*2048+1179,   37*2048+1180,    5*2048+1181,   11*2048+1182,   45*2048+1183,   43*2048+1184,   36*2048+1185,   45*2048+1186,   45*2048+1187, 
  16*2048+1188,   43*2048+1189,    1*2048+1190,   24*2048+1191,   19*2048+1192,   28*2048+1193,   45*2048+1194,   30*2048+1195,   11*2048+1196,   45*2048+1197,   45*2048+1198, 
  35*2048+1199,   11*2048+1200,    5*2048+1201,   17*2048+1202,   30*2048+1203,   45*2048+1204,   16*2048+1205,    0*2048+1206,   31*2048+1207,   45*2048+1208,   45*2048+1209, 
  43*2048+1210,   39*2048+1211,   14*2048+1212,   34*2048+1213,    6*2048+1214,   39*2048+1215,   45*2048+1216,    1*2048+1217,   17*2048+1218,   45*2048+1219,   45*2048+1220, 
  38*2048+1221,   24*2048+1222,   16*2048+1223,   35*2048+1224,   40*2048+1225,    2*2048+1226,   45*2048+1227,    6*2048+1228,    4*2048+1229,   45*2048+1230,   45*2048+1231, 
  42*2048+1232,   37*2048+1233,   26*2048+1234,    6*2048+1235,   22*2048+1236,   33*2048+1237,   30*2048+1238,   45*2048+1239,   12*2048+1240,   45*2048+1241,   45*2048+1242, 
  38*2048+1243,   12*2048+1244,   45*2048+1245,   27*2048+1246,   25*2048+1247,   12*2048+1248,   45*2048+1249,   33*2048+1250,   41*2048+1251,   45*2048+1252,   45*2048+1253, 
   9*2048+1254,   36*2048+1255,   27*2048+1256,   36*2048+1257,   15*2048+1258,   19*2048+1259,   30*2048+1260,    9*2048+1261,   45*2048+1262,   45*2048+1263,   45*2048+1264, 
   6*2048+1265,   40*2048+1266,   23*2048+1267,   27*2048+1268,   11*2048+1269,   16*2048+1270,   29*2048+1271,   45*2048+1272,   23*2048+1273,   45*2048+1274,   45*2048+1275, 
  16*2048+1276,   19*2048+1277,    7*2048+1278,   25*2048+1279,    6*2048+1280,   45*2048+1281,   15*2048+1282,   11*2048+1283,   20*2048+1284,   45*2048+1285,   45*2048+1286, 
  25*2048+1287,   23*2048+1288,   10*2048+1289,   13*2048+1290,    8*2048+1291,    4*2048+1292,   19*2048+1293,   45*2048+1294,   16*2048+1295,   45*2048+1296,   45*2048+1297, 
   4*2048+1298,   28*2048+1299,   22*2048+1300,   22*2048+1301,   32*2048+1302,    2*2048+1303,   14*2048+1304,   45*2048+1305,   19*2048+1306,   45*2048+1307,   45*2048+1308, 
  18*2048+1309,   31*2048+1310,   26*2048+1311,   29*2048+1312,   39*2048+1313,   45*2048+1314,   12*2048+1315,   28*2048+1316,   33*2048+1317,   45*2048+1318,   45*2048+1319, 
  33*2048+1320,   36*2048+1321,   44*2048+1322,   30*2048+1323,   25*2048+1324,    6*2048+1325,    1*2048+1326,   45*2048+1327,   11*2048+1328,   45*2048+1329,   45*2048+1330, 
  44*2048+1331,   34*2048+1332,   44*2048+1333,    5*2048+1334,   38*2048+1335,   18*2048+1336,   18*2048+1337,   45*2048+1338,   20*2048+1339,   45*2048+1340,   45*2048+1341, 
  13*2048+1342,   44*2048+1343,   26*2048+1344,   18*2048+1345,   16*2048+1346,    3*2048+1347,   45*2048+1348,   20*2048+1349,   42*2048+1350,   45*2048+1351,   45*2048+1352, 
   6*2048+1353,   37*2048+1354,   22*2048+1355,   21*2048+1356,    8*2048+1357,   10*2048+1358,   40*2048+1359,   45*2048+1360,    3*2048+1361,   45*2048+1362,   45*2048+1363, 
  29*2048+1364,   13*2048+1365,    4*2048+1366,   16*2048+1367,   14*2048+1368,   18*2048+1369,   40*2048+1370,   45*2048+1371,    1*2048+1372,   45*2048+1373,   45*2048+1374, 
  20*2048+1375,    4*2048+1376,   25*2048+1377,   37*2048+1378,    5*2048+1379,   11*2048+1380,   45*2048+1381,   43*2048+1382,   36*2048+1383,   45*2048+1384,   45*2048+1385, 
  31*2048+1386,   12*2048+1387,   16*2048+1388,   43*2048+1389,    1*2048+1390,   24*2048+1391,   19*2048+1392,   28*2048+1393,   45*2048+1394,   45*2048+1395,   45*2048+1396, 
   1*2048+1397,   32*2048+1398,   35*2048+1399,   11*2048+1400,    5*2048+1401,   17*2048+1402,   30*2048+1403,   45*2048+1404,   16*2048+1405,   45*2048+1406,   45*2048+1407, 
   2*2048+1408,   18*2048+1409,   43*2048+1410,   39*2048+1411,   14*2048+1412,   34*2048+1413,    6*2048+1414,   39*2048+1415,   45*2048+1416,   45*2048+1417,   45*2048+1418, 
   7*2048+1419,    5*2048+1420,   38*2048+1421,   24*2048+1422,   16*2048+1423,   35*2048+1424,   40*2048+1425,    2*2048+1426,   45*2048+1427,   45*2048+1428,   45*2048+1429, 
  13*2048+1430,   42*2048+1431,   37*2048+1432,   26*2048+1433,    6*2048+1434,   22*2048+1435,   33*2048+1436,   30*2048+1437,   45*2048+1438,   45*2048+1439,   45*2048+1440, 
  42*2048+1441,   38*2048+1442,   12*2048+1443,   45*2048+1444,   27*2048+1445,   25*2048+1446,   12*2048+1447,   45*2048+1448,   33*2048+1449,   45*2048+1450,   45*2048+1451, 
   9*2048+1452,   36*2048+1453,   27*2048+1454,   36*2048+1455,   15*2048+1456,   19*2048+1457,   30*2048+1458,    9*2048+1459,   45*2048+1460,   45*2048+1461,   45*2048+1462, 
  24*2048+1463,    6*2048+1464,   40*2048+1465,   23*2048+1466,   27*2048+1467,   11*2048+1468,   16*2048+1469,   29*2048+1470,   45*2048+1471,   45*2048+1472,   45*2048+1473, 
  16*2048+1474,   12*2048+1475,   21*2048+1476,   16*2048+1477,   19*2048+1478,    7*2048+1479,   25*2048+1480,    6*2048+1481,   45*2048+1482,   45*2048+1483,   45*2048+1484, 
  17*2048+1485,   25*2048+1486,   23*2048+1487,   10*2048+1488,   13*2048+1489,    8*2048+1490,    4*2048+1491,   19*2048+1492,   45*2048+1493,   45*2048+1494,   45*2048+1495, 
  20*2048+1496,    4*2048+1497,   28*2048+1498,   22*2048+1499,   22*2048+1500,   32*2048+1501,    2*2048+1502,   14*2048+1503,   45*2048+1504,   45*2048+1505,   45*2048+1506, 
  29*2048+1507,   34*2048+1508,   18*2048+1509,   31*2048+1510,   26*2048+1511,   29*2048+1512,   39*2048+1513,   45*2048+1514,   12*2048+1515,   45*2048+1516,   45*2048+1517, 
  33*2048+1518,   36*2048+1519,   44*2048+1520,   30*2048+1521,   25*2048+1522,    6*2048+1523,    1*2048+1524,   45*2048+1525,   11*2048+1526,   45*2048+1527,   45*2048+1528, 
  21*2048+1529,   44*2048+1530,   34*2048+1531,   44*2048+1532,    5*2048+1533,   38*2048+1534,   18*2048+1535,   18*2048+1536,   45*2048+1537,   45*2048+1538,   45*2048+1539, 
  21*2048+1540,   43*2048+1541,   13*2048+1542,   44*2048+1543,   26*2048+1544,   18*2048+1545,   16*2048+1546,    3*2048+1547,   45*2048+1548,   45*2048+1549,   45*2048+1550, 
   4*2048+1551,    6*2048+1552,   37*2048+1553,   22*2048+1554,   21*2048+1555,    8*2048+1556,   10*2048+1557,   40*2048+1558,   45*2048+1559,   45*2048+1560,   45*2048+1561, 
   2*2048+1562,   29*2048+1563,   13*2048+1564,    4*2048+1565,   16*2048+1566,   14*2048+1567,   18*2048+1568,   40*2048+1569,   45*2048+1570,   45*2048+1571,   45*2048+1572, 
  44*2048+1573,   37*2048+1574,   20*2048+1575,    4*2048+1576,   25*2048+1577,   37*2048+1578,    5*2048+1579,   11*2048+1580,   45*2048+1581,   45*2048+1582,   45*2048+1583, 

  45*2048+   0,   21*2048+   1,   45*2048+   2,   32*2048+   3,   39*2048+   4,   21*2048+   5,    6*2048+   6,   36*2048+   7,   45*2048+   8,   44*2048+   9, 
  45*2048+  10,   45*2048+  11,   43*2048+  12,   16*2048+  13,   18*2048+  14,   32*2048+  15,    6*2048+  16,   23*2048+  17,   45*2048+  18,   45*2048+  19, 
  44*2048+  20,   45*2048+  21,   45*2048+  22,   44*2048+  23,   27*2048+  24,   42*2048+  25,    2*2048+  26,   29*2048+  27,   45*2048+  28,   45*2048+  29, 
  45*2048+  30,   43*2048+  31,   45*2048+  32,   32*2048+  33,   19*2048+  34,   30*2048+  35,   23*2048+  36,   20*2048+  37,   45*2048+  38,   45*2048+  39, 
  45*2048+  40,   45*2048+  41,   31*2048+  42,   13*2048+  43,   15*2048+  44,   15*2048+  45,   35*2048+  46,   42*2048+  47,   45*2048+  48,   45*2048+  49, 
  19*2048+  50,   45*2048+  51,   45*2048+  52,    4*2048+  53,   29*2048+  54,   31*2048+  55,   39*2048+  56,   32*2048+  57,   45*2048+  58,   45*2048+  59, 
  45*2048+  60,   45*2048+  61,   43*2048+  62,    9*2048+  63,   24*2048+  64,   16*2048+  65,   11*2048+  66,    4*2048+  67,   45*2048+  68,   45*2048+  69, 
   1*2048+  70,   45*2048+  71,   27*2048+  72,   45*2048+  73,   41*2048+  74,   24*2048+  75,    9*2048+  76,    1*2048+  77,   45*2048+  78,   45*2048+  79, 
  45*2048+  80,   13*2048+  81,   45*2048+  82,   13*2048+  83,    8*2048+  84,   40*2048+  85,   31*2048+  86,    8*2048+  87,   45*2048+  88,   45*2048+  89, 
  17*2048+  90,   45*2048+  91,   45*2048+  92,   25*2048+  93,   12*2048+  94,   16*2048+  95,   37*2048+  96,   12*2048+  97,   45*2048+  98,   45*2048+  99, 
  23*2048+ 100,   45*2048+ 101,   45*2048+ 102,   27*2048+ 103,   35*2048+ 104,   25*2048+ 105,   25*2048+ 106,   33*2048+ 107,   45*2048+ 108,   45*2048+ 109, 
  37*2048+ 110,   20*2048+ 111,   45*2048+ 112,   45*2048+ 113,   33*2048+ 114,   34*2048+ 115,   12*2048+ 116,   22*2048+ 117,   45*2048+ 118,   45*2048+ 119, 
  45*2048+ 120,   45*2048+ 121,   23*2048+ 122,   42*2048+ 123,   32*2048+ 124,   32*2048+ 125,   33*2048+ 126,   20*2048+ 127,   45*2048+ 128,   45*2048+ 129, 
  42*2048+ 130,   45*2048+ 131,   45*2048+ 132,   10*2048+ 133,   16*2048+ 134,   39*2048+ 135,   36*2048+ 136,   43*2048+ 137,   45*2048+ 138,   45*2048+ 139, 
  45*2048+ 140,   45*2048+ 141,   37*2048+ 142,   24*2048+ 143,   27*2048+ 144,   43*2048+ 145,   40*2048+ 146,   43*2048+ 147,   45*2048+ 148,   45*2048+ 149, 
  45*2048+ 150,   21*2048+ 151,   45*2048+ 152,   32*2048+ 153,   39*2048+ 154,   21*2048+ 155,    6*2048+ 156,   36*2048+ 157,   45*2048+ 158,   45*2048+ 159, 
  24*2048+ 160,   45*2048+ 161,   45*2048+ 162,   43*2048+ 163,   16*2048+ 164,   18*2048+ 165,   32*2048+ 166,    6*2048+ 167,   45*2048+ 168,   45*2048+ 169, 
  44*2048+ 170,   45*2048+ 171,   45*2048+ 172,   44*2048+ 173,   27*2048+ 174,   42*2048+ 175,    2*2048+ 176,   29*2048+ 177,   45*2048+ 178,   45*2048+ 179, 
  45*2048+ 180,   43*2048+ 181,   45*2048+ 182,   32*2048+ 183,   19*2048+ 184,   30*2048+ 185,   23*2048+ 186,   20*2048+ 187,   45*2048+ 188,   45*2048+ 189, 
  43*2048+ 190,   45*2048+ 191,   45*2048+ 192,   31*2048+ 193,   13*2048+ 194,   15*2048+ 195,   15*2048+ 196,   35*2048+ 197,   45*2048+ 198,   45*2048+ 199, 
  33*2048+ 200,   19*2048+ 201,   45*2048+ 202,   45*2048+ 203,    4*2048+ 204,   29*2048+ 205,   31*2048+ 206,   39*2048+ 207,   45*2048+ 208,   45*2048+ 209, 
  45*2048+ 210,   45*2048+ 211,   43*2048+ 212,    9*2048+ 213,   24*2048+ 214,   16*2048+ 215,   11*2048+ 216,    4*2048+ 217,   45*2048+ 218,   45*2048+ 219, 
   1*2048+ 220,   45*2048+ 221,   27*2048+ 222,   45*2048+ 223,   41*2048+ 224,   24*2048+ 225,    9*2048+ 226,    1*2048+ 227,   45*2048+ 228,   45*2048+ 229, 
  45*2048+ 230,   13*2048+ 231,   45*2048+ 232,   13*2048+ 233,    8*2048+ 234,   40*2048+ 235,   31*2048+ 236,    8*2048+ 237,   45*2048+ 238,   45*2048+ 239, 
  38*2048+ 240,   13*2048+ 241,   17*2048+ 242,   45*2048+ 243,   45*2048+ 244,   25*2048+ 245,   12*2048+ 246,   16*2048+ 247,   45*2048+ 248,   45*2048+ 249, 
  23*2048+ 250,   45*2048+ 251,   45*2048+ 252,   27*2048+ 253,   35*2048+ 254,   25*2048+ 255,   25*2048+ 256,   33*2048+ 257,   45*2048+ 258,   45*2048+ 259, 
  37*2048+ 260,   20*2048+ 261,   45*2048+ 262,   45*2048+ 263,   33*2048+ 264,   34*2048+ 265,   12*2048+ 266,   22*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
  45*2048+ 270,   45*2048+ 271,   23*2048+ 272,   42*2048+ 273,   32*2048+ 274,   32*2048+ 275,   33*2048+ 276,   20*2048+ 277,   45*2048+ 278,   45*2048+ 279, 
  42*2048+ 280,   45*2048+ 281,   45*2048+ 282,   10*2048+ 283,   16*2048+ 284,   39*2048+ 285,   36*2048+ 286,   43*2048+ 287,   45*2048+ 288,   45*2048+ 289, 
  41*2048+ 290,   44*2048+ 291,   45*2048+ 292,   45*2048+ 293,   37*2048+ 294,   24*2048+ 295,   27*2048+ 296,   43*2048+ 297,   45*2048+ 298,   45*2048+ 299, 
  45*2048+ 300,   21*2048+ 301,   45*2048+ 302,   32*2048+ 303,   39*2048+ 304,   21*2048+ 305,    6*2048+ 306,   36*2048+ 307,   45*2048+ 308,   45*2048+ 309, 
  24*2048+ 310,   45*2048+ 311,   45*2048+ 312,   43*2048+ 313,   16*2048+ 314,   18*2048+ 315,   32*2048+ 316,    6*2048+ 317,   45*2048+ 318,   45*2048+ 319, 
  44*2048+ 320,   45*2048+ 321,   45*2048+ 322,   44*2048+ 323,   27*2048+ 324,   42*2048+ 325,    2*2048+ 326,   29*2048+ 327,   45*2048+ 328,   45*2048+ 329, 
  45*2048+ 330,   43*2048+ 331,   45*2048+ 332,   32*2048+ 333,   19*2048+ 334,   30*2048+ 335,   23*2048+ 336,   20*2048+ 337,   45*2048+ 338,   45*2048+ 339, 
  43*2048+ 340,   45*2048+ 341,   45*2048+ 342,   31*2048+ 343,   13*2048+ 344,   15*2048+ 345,   15*2048+ 346,   35*2048+ 347,   45*2048+ 348,   45*2048+ 349, 
  40*2048+ 350,   33*2048+ 351,   19*2048+ 352,   45*2048+ 353,   45*2048+ 354,    4*2048+ 355,   29*2048+ 356,   31*2048+ 357,   45*2048+ 358,   45*2048+ 359, 
  12*2048+ 360,    5*2048+ 361,   45*2048+ 362,   45*2048+ 363,   43*2048+ 364,    9*2048+ 365,   24*2048+ 366,   16*2048+ 367,   45*2048+ 368,   45*2048+ 369, 
   1*2048+ 370,   45*2048+ 371,   27*2048+ 372,   45*2048+ 373,   41*2048+ 374,   24*2048+ 375,    9*2048+ 376,    1*2048+ 377,   45*2048+ 378,   45*2048+ 379, 
   9*2048+ 380,   45*2048+ 381,   13*2048+ 382,   45*2048+ 383,   13*2048+ 384,    8*2048+ 385,   40*2048+ 386,   31*2048+ 387,   45*2048+ 388,   45*2048+ 389, 
  17*2048+ 390,   38*2048+ 391,   13*2048+ 392,   17*2048+ 393,   45*2048+ 394,   45*2048+ 395,   25*2048+ 396,   12*2048+ 397,   45*2048+ 398,   45*2048+ 399, 
  34*2048+ 400,   23*2048+ 401,   45*2048+ 402,   45*2048+ 403,   27*2048+ 404,   35*2048+ 405,   25*2048+ 406,   25*2048+ 407,   45*2048+ 408,   45*2048+ 409, 
  37*2048+ 410,   20*2048+ 411,   45*2048+ 412,   45*2048+ 413,   33*2048+ 414,   34*2048+ 415,   12*2048+ 416,   22*2048+ 417,   45*2048+ 418,   45*2048+ 419, 
  21*2048+ 420,   45*2048+ 421,   45*2048+ 422,   23*2048+ 423,   42*2048+ 424,   32*2048+ 425,   32*2048+ 426,   33*2048+ 427,   45*2048+ 428,   45*2048+ 429, 
  37*2048+ 430,   44*2048+ 431,   42*2048+ 432,   45*2048+ 433,   45*2048+ 434,   10*2048+ 435,   16*2048+ 436,   39*2048+ 437,   45*2048+ 438,   45*2048+ 439, 
  28*2048+ 440,   44*2048+ 441,   41*2048+ 442,   44*2048+ 443,   45*2048+ 444,   45*2048+ 445,   37*2048+ 446,   24*2048+ 447,   45*2048+ 448,   45*2048+ 449, 
  37*2048+ 450,   45*2048+ 451,   21*2048+ 452,   45*2048+ 453,   32*2048+ 454,   39*2048+ 455,   21*2048+ 456,    6*2048+ 457,   45*2048+ 458,   45*2048+ 459, 
   7*2048+ 460,   24*2048+ 461,   45*2048+ 462,   45*2048+ 463,   43*2048+ 464,   16*2048+ 465,   18*2048+ 466,   32*2048+ 467,   45*2048+ 468,   45*2048+ 469, 
  30*2048+ 470,   44*2048+ 471,   45*2048+ 472,   45*2048+ 473,   44*2048+ 474,   27*2048+ 475,   42*2048+ 476,    2*2048+ 477,   45*2048+ 478,   45*2048+ 479, 
  21*2048+ 480,   45*2048+ 481,   43*2048+ 482,   45*2048+ 483,   32*2048+ 484,   19*2048+ 485,   30*2048+ 486,   23*2048+ 487,   45*2048+ 488,   45*2048+ 489, 
  16*2048+ 490,   16*2048+ 491,   36*2048+ 492,   43*2048+ 493,   45*2048+ 494,   45*2048+ 495,   31*2048+ 496,   13*2048+ 497,   45*2048+ 498,   45*2048+ 499, 
  40*2048+ 500,   33*2048+ 501,   19*2048+ 502,   45*2048+ 503,   45*2048+ 504,    4*2048+ 505,   29*2048+ 506,   31*2048+ 507,   45*2048+ 508,   45*2048+ 509, 
  12*2048+ 510,    5*2048+ 511,   45*2048+ 512,   45*2048+ 513,   43*2048+ 514,    9*2048+ 515,   24*2048+ 516,   16*2048+ 517,   45*2048+ 518,   45*2048+ 519, 
   2*2048+ 520,    1*2048+ 521,   45*2048+ 522,   27*2048+ 523,   45*2048+ 524,   41*2048+ 525,   24*2048+ 526,    9*2048+ 527,   45*2048+ 528,   45*2048+ 529, 
  32*2048+ 530,    9*2048+ 531,   45*2048+ 532,   13*2048+ 533,   45*2048+ 534,   13*2048+ 535,    8*2048+ 536,   40*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
  13*2048+ 540,   17*2048+ 541,   38*2048+ 542,   13*2048+ 543,   17*2048+ 544,   45*2048+ 545,   45*2048+ 546,   25*2048+ 547,   45*2048+ 548,   45*2048+ 549, 
  34*2048+ 550,   23*2048+ 551,   45*2048+ 552,   45*2048+ 553,   27*2048+ 554,   35*2048+ 555,   25*2048+ 556,   25*2048+ 557,   45*2048+ 558,   45*2048+ 559, 
  23*2048+ 560,   37*2048+ 561,   20*2048+ 562,   45*2048+ 563,   45*2048+ 564,   33*2048+ 565,   34*2048+ 566,   12*2048+ 567,   45*2048+ 568,   45*2048+ 569, 
  21*2048+ 570,   45*2048+ 571,   45*2048+ 572,   23*2048+ 573,   42*2048+ 574,   32*2048+ 575,   32*2048+ 576,   33*2048+ 577,   45*2048+ 578,   45*2048+ 579, 
  37*2048+ 580,   44*2048+ 581,   42*2048+ 582,   45*2048+ 583,   45*2048+ 584,   10*2048+ 585,   16*2048+ 586,   39*2048+ 587,   45*2048+ 588,   45*2048+ 589, 
  28*2048+ 590,   44*2048+ 591,   41*2048+ 592,   44*2048+ 593,   45*2048+ 594,   45*2048+ 595,   37*2048+ 596,   24*2048+ 597,   45*2048+ 598,   45*2048+ 599, 
   7*2048+ 600,   37*2048+ 601,   45*2048+ 602,   21*2048+ 603,   45*2048+ 604,   32*2048+ 605,   39*2048+ 606,   21*2048+ 607,   45*2048+ 608,   45*2048+ 609, 
   7*2048+ 610,   24*2048+ 611,   45*2048+ 612,   45*2048+ 613,   43*2048+ 614,   16*2048+ 615,   18*2048+ 616,   32*2048+ 617,   45*2048+ 618,   45*2048+ 619, 
  30*2048+ 620,   44*2048+ 621,   45*2048+ 622,   45*2048+ 623,   44*2048+ 624,   27*2048+ 625,   42*2048+ 626,    2*2048+ 627,   45*2048+ 628,   45*2048+ 629, 
  31*2048+ 630,   24*2048+ 631,   21*2048+ 632,   45*2048+ 633,   43*2048+ 634,   45*2048+ 635,   32*2048+ 636,   19*2048+ 637,   45*2048+ 638,   45*2048+ 639, 
  16*2048+ 640,   16*2048+ 641,   36*2048+ 642,   43*2048+ 643,   45*2048+ 644,   45*2048+ 645,   31*2048+ 646,   13*2048+ 647,   45*2048+ 648,   45*2048+ 649, 
  40*2048+ 650,   33*2048+ 651,   19*2048+ 652,   45*2048+ 653,   45*2048+ 654,    4*2048+ 655,   29*2048+ 656,   31*2048+ 657,   45*2048+ 658,   45*2048+ 659, 
  17*2048+ 660,   12*2048+ 661,    5*2048+ 662,   45*2048+ 663,   45*2048+ 664,   43*2048+ 665,    9*2048+ 666,   24*2048+ 667,   45*2048+ 668,   45*2048+ 669, 
   2*2048+ 670,    1*2048+ 671,   45*2048+ 672,   27*2048+ 673,   45*2048+ 674,   41*2048+ 675,   24*2048+ 676,    9*2048+ 677,   45*2048+ 678,   45*2048+ 679, 
  32*2048+ 680,    9*2048+ 681,   45*2048+ 682,   13*2048+ 683,   45*2048+ 684,   13*2048+ 685,    8*2048+ 686,   40*2048+ 687,   45*2048+ 688,   45*2048+ 689, 
  13*2048+ 690,   17*2048+ 691,   38*2048+ 692,   13*2048+ 693,   17*2048+ 694,   45*2048+ 695,   45*2048+ 696,   25*2048+ 697,   45*2048+ 698,   45*2048+ 699, 
  26*2048+ 700,   34*2048+ 701,   23*2048+ 702,   45*2048+ 703,   45*2048+ 704,   27*2048+ 705,   35*2048+ 706,   25*2048+ 707,   45*2048+ 708,   45*2048+ 709, 
  23*2048+ 710,   37*2048+ 711,   20*2048+ 712,   45*2048+ 713,   45*2048+ 714,   33*2048+ 715,   34*2048+ 716,   12*2048+ 717,   45*2048+ 718,   45*2048+ 719, 
  21*2048+ 720,   45*2048+ 721,   45*2048+ 722,   23*2048+ 723,   42*2048+ 724,   32*2048+ 725,   32*2048+ 726,   33*2048+ 727,   45*2048+ 728,   45*2048+ 729, 
  37*2048+ 730,   44*2048+ 731,   42*2048+ 732,   45*2048+ 733,   45*2048+ 734,   10*2048+ 735,   16*2048+ 736,   39*2048+ 737,   45*2048+ 738,   45*2048+ 739, 
  25*2048+ 740,   28*2048+ 741,   44*2048+ 742,   41*2048+ 743,   44*2048+ 744,   45*2048+ 745,   45*2048+ 746,   37*2048+ 747,   45*2048+ 748,   45*2048+ 749, 
  22*2048+ 750,    7*2048+ 751,   37*2048+ 752,   45*2048+ 753,   21*2048+ 754,   45*2048+ 755,   32*2048+ 756,   39*2048+ 757,   45*2048+ 758,   45*2048+ 759, 
  19*2048+ 760,   33*2048+ 761,    7*2048+ 762,   24*2048+ 763,   45*2048+ 764,   45*2048+ 765,   43*2048+ 766,   16*2048+ 767,   45*2048+ 768,   45*2048+ 769, 
   3*2048+ 770,   30*2048+ 771,   44*2048+ 772,   45*2048+ 773,   45*2048+ 774,   44*2048+ 775,   27*2048+ 776,   42*2048+ 777,   45*2048+ 778,   45*2048+ 779, 
  31*2048+ 780,   24*2048+ 781,   21*2048+ 782,   45*2048+ 783,   43*2048+ 784,   45*2048+ 785,   32*2048+ 786,   19*2048+ 787,   45*2048+ 788,   45*2048+ 789, 
  14*2048+ 790,   16*2048+ 791,   16*2048+ 792,   36*2048+ 793,   43*2048+ 794,   45*2048+ 795,   45*2048+ 796,   31*2048+ 797,   45*2048+ 798,   45*2048+ 799, 
  30*2048+ 800,   32*2048+ 801,   40*2048+ 802,   33*2048+ 803,   19*2048+ 804,   45*2048+ 805,   45*2048+ 806,    4*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  25*2048+ 810,   17*2048+ 811,   12*2048+ 812,    5*2048+ 813,   45*2048+ 814,   45*2048+ 815,   43*2048+ 816,    9*2048+ 817,   45*2048+ 818,   45*2048+ 819, 
   2*2048+ 820,    1*2048+ 821,   45*2048+ 822,   27*2048+ 823,   45*2048+ 824,   41*2048+ 825,   24*2048+ 826,    9*2048+ 827,   45*2048+ 828,   45*2048+ 829, 
  41*2048+ 830,   32*2048+ 831,    9*2048+ 832,   45*2048+ 833,   13*2048+ 834,   45*2048+ 835,   13*2048+ 836,    8*2048+ 837,   45*2048+ 838,   45*2048+ 839, 
  26*2048+ 840,   13*2048+ 841,   17*2048+ 842,   38*2048+ 843,   13*2048+ 844,   17*2048+ 845,   45*2048+ 846,   45*2048+ 847,   45*2048+ 848,   45*2048+ 849, 
  26*2048+ 850,   26*2048+ 851,   34*2048+ 852,   23*2048+ 853,   45*2048+ 854,   45*2048+ 855,   27*2048+ 856,   35*2048+ 857,   45*2048+ 858,   45*2048+ 859, 
  35*2048+ 860,   13*2048+ 861,   23*2048+ 862,   37*2048+ 863,   20*2048+ 864,   45*2048+ 865,   45*2048+ 866,   33*2048+ 867,   45*2048+ 868,   45*2048+ 869, 
  34*2048+ 870,   21*2048+ 871,   45*2048+ 872,   45*2048+ 873,   23*2048+ 874,   42*2048+ 875,   32*2048+ 876,   32*2048+ 877,   45*2048+ 878,   45*2048+ 879, 
  17*2048+ 880,   40*2048+ 881,   37*2048+ 882,   44*2048+ 883,   42*2048+ 884,   45*2048+ 885,   45*2048+ 886,   10*2048+ 887,   45*2048+ 888,   45*2048+ 889, 
  38*2048+ 890,   25*2048+ 891,   28*2048+ 892,   44*2048+ 893,   41*2048+ 894,   44*2048+ 895,   45*2048+ 896,   45*2048+ 897,   45*2048+ 898,   45*2048+ 899, 
  22*2048+ 900,    7*2048+ 901,   37*2048+ 902,   45*2048+ 903,   21*2048+ 904,   45*2048+ 905,   32*2048+ 906,   39*2048+ 907,   45*2048+ 908,   45*2048+ 909, 
  17*2048+ 910,   19*2048+ 911,   33*2048+ 912,    7*2048+ 913,   24*2048+ 914,   45*2048+ 915,   45*2048+ 916,   43*2048+ 917,   45*2048+ 918,   45*2048+ 919, 
   3*2048+ 920,   30*2048+ 921,   44*2048+ 922,   45*2048+ 923,   45*2048+ 924,   44*2048+ 925,   27*2048+ 926,   42*2048+ 927,   45*2048+ 928,   45*2048+ 929, 
  31*2048+ 930,   24*2048+ 931,   21*2048+ 932,   45*2048+ 933,   43*2048+ 934,   45*2048+ 935,   32*2048+ 936,   19*2048+ 937,   45*2048+ 938,   45*2048+ 939, 
  14*2048+ 940,   16*2048+ 941,   16*2048+ 942,   36*2048+ 943,   43*2048+ 944,   45*2048+ 945,   45*2048+ 946,   31*2048+ 947,   45*2048+ 948,   45*2048+ 949, 
  30*2048+ 950,   32*2048+ 951,   40*2048+ 952,   33*2048+ 953,   19*2048+ 954,   45*2048+ 955,   45*2048+ 956,    4*2048+ 957,   45*2048+ 958,   45*2048+ 959, 
  10*2048+ 960,   25*2048+ 961,   17*2048+ 962,   12*2048+ 963,    5*2048+ 964,   45*2048+ 965,   45*2048+ 966,   43*2048+ 967,   45*2048+ 968,   45*2048+ 969, 
  10*2048+ 970,    2*2048+ 971,    1*2048+ 972,   45*2048+ 973,   27*2048+ 974,   45*2048+ 975,   41*2048+ 976,   24*2048+ 977,   45*2048+ 978,   45*2048+ 979, 
   9*2048+ 980,   41*2048+ 981,   32*2048+ 982,    9*2048+ 983,   45*2048+ 984,   13*2048+ 985,   45*2048+ 986,   13*2048+ 987,   45*2048+ 988,   45*2048+ 989, 
  26*2048+ 990,   13*2048+ 991,   17*2048+ 992,   38*2048+ 993,   13*2048+ 994,   17*2048+ 995,   45*2048+ 996,   45*2048+ 997,   45*2048+ 998,   45*2048+ 999, 
  36*2048+1000,   26*2048+1001,   26*2048+1002,   34*2048+1003,   23*2048+1004,   45*2048+1005,   45*2048+1006,   27*2048+1007,   45*2048+1008,   45*2048+1009, 
  35*2048+1010,   13*2048+1011,   23*2048+1012,   37*2048+1013,   20*2048+1014,   45*2048+1015,   45*2048+1016,   33*2048+1017,   45*2048+1018,   45*2048+1019, 
  24*2048+1020,   43*2048+1021,   33*2048+1022,   33*2048+1023,   34*2048+1024,   21*2048+1025,   45*2048+1026,   45*2048+1027,   45*2048+1028,   45*2048+1029, 
  17*2048+1030,   40*2048+1031,   37*2048+1032,   44*2048+1033,   42*2048+1034,   45*2048+1035,   45*2048+1036,   10*2048+1037,   45*2048+1038,   45*2048+1039, 
  38*2048+1040,   25*2048+1041,   28*2048+1042,   44*2048+1043,   41*2048+1044,   44*2048+1045,   45*2048+1046,   45*2048+1047,   45*2048+1048,   45*2048+1049, 
  40*2048+1050,   22*2048+1051,    7*2048+1052,   37*2048+1053,   45*2048+1054,   21*2048+1055,   45*2048+1056,   32*2048+1057,   45*2048+1058,   45*2048+1059, 
  44*2048+1060,   17*2048+1061,   19*2048+1062,   33*2048+1063,    7*2048+1064,   24*2048+1065,   45*2048+1066,   45*2048+1067,   45*2048+1068,   45*2048+1069, 
  45*2048+1070,   28*2048+1071,   43*2048+1072,    3*2048+1073,   30*2048+1074,   44*2048+1075,   45*2048+1076,   45*2048+1077,   45*2048+1078,   45*2048+1079, 
  33*2048+1080,   20*2048+1081,   31*2048+1082,   24*2048+1083,   21*2048+1084,   45*2048+1085,   43*2048+1086,   45*2048+1087,   45*2048+1088,   45*2048+1089, 
  14*2048+1090,   16*2048+1091,   16*2048+1092,   36*2048+1093,   43*2048+1094,   45*2048+1095,   45*2048+1096,   31*2048+1097,   45*2048+1098,   45*2048+1099, 
   5*2048+1100,   30*2048+1101,   32*2048+1102,   40*2048+1103,   33*2048+1104,   19*2048+1105,   45*2048+1106,   45*2048+1107,   45*2048+1108,   45*2048+1109, 
  44*2048+1110,   10*2048+1111,   25*2048+1112,   17*2048+1113,   12*2048+1114,    5*2048+1115,   45*2048+1116,   45*2048+1117,   45*2048+1118,   45*2048+1119, 
  25*2048+1120,   10*2048+1121,    2*2048+1122,    1*2048+1123,   45*2048+1124,   27*2048+1125,   45*2048+1126,   41*2048+1127,   45*2048+1128,   45*2048+1129, 
  14*2048+1130,    9*2048+1131,   41*2048+1132,   32*2048+1133,    9*2048+1134,   45*2048+1135,   13*2048+1136,   45*2048+1137,   45*2048+1138,   45*2048+1139, 
  26*2048+1140,   13*2048+1141,   17*2048+1142,   38*2048+1143,   13*2048+1144,   17*2048+1145,   45*2048+1146,   45*2048+1147,   45*2048+1148,   45*2048+1149, 
  28*2048+1150,   36*2048+1151,   26*2048+1152,   26*2048+1153,   34*2048+1154,   23*2048+1155,   45*2048+1156,   45*2048+1157,   45*2048+1158,   45*2048+1159, 
  34*2048+1160,   35*2048+1161,   13*2048+1162,   23*2048+1163,   37*2048+1164,   20*2048+1165,   45*2048+1166,   45*2048+1167,   45*2048+1168,   45*2048+1169, 
  24*2048+1170,   43*2048+1171,   33*2048+1172,   33*2048+1173,   34*2048+1174,   21*2048+1175,   45*2048+1176,   45*2048+1177,   45*2048+1178,   45*2048+1179, 
  11*2048+1180,   17*2048+1181,   40*2048+1182,   37*2048+1183,   44*2048+1184,   42*2048+1185,   45*2048+1186,   45*2048+1187,   45*2048+1188,   45*2048+1189, 
  38*2048+1190,   25*2048+1191,   28*2048+1192,   44*2048+1193,   41*2048+1194,   44*2048+1195,   45*2048+1196,   45*2048+1197,   45*2048+1198,   45*2048+1199, 

  45*2048+  33,   45*2048+  34,   45*2048+  35,    9*2048+  36,    4*2048+  37,   38*2048+  38,   13*2048+  39,   45*2048+  40,   45*2048+  41, 
  45*2048+ 165,   45*2048+ 166,   45*2048+ 167,    9*2048+ 168,    4*2048+ 169,   38*2048+ 170,   13*2048+ 171,   45*2048+ 172,   45*2048+ 173, 
  14*2048+ 297,   45*2048+ 298,   45*2048+ 299,   45*2048+ 300,    9*2048+ 301,    4*2048+ 302,   38*2048+ 303,   45*2048+ 304,   45*2048+ 305, 
  39*2048+ 429,   14*2048+ 430,   45*2048+ 431,   45*2048+ 432,   45*2048+ 433,    9*2048+ 434,    4*2048+ 435,   45*2048+ 436,   45*2048+ 437, 
  39*2048+ 561,   14*2048+ 562,   45*2048+ 563,   45*2048+ 564,   45*2048+ 565,    9*2048+ 566,    4*2048+ 567,   45*2048+ 568,   45*2048+ 569, 
   5*2048+ 693,   39*2048+ 694,   14*2048+ 695,   45*2048+ 696,   45*2048+ 697,   45*2048+ 698,    9*2048+ 699,   45*2048+ 700,   45*2048+ 701, 
   5*2048+ 825,   39*2048+ 826,   14*2048+ 827,   45*2048+ 828,   45*2048+ 829,   45*2048+ 830,    9*2048+ 831,   45*2048+ 832,   45*2048+ 833, 
  10*2048+ 957,    5*2048+ 958,   39*2048+ 959,   14*2048+ 960,   45*2048+ 961,   45*2048+ 962,   45*2048+ 963,   45*2048+ 964,   45*2048+ 965, 
  45*2048+   0,   45*2048+   1,   27*2048+   2,   43*2048+   3,   18*2048+   4,   17*2048+   5,   34*2048+   6,   15*2048+   7,   45*2048+   8,   44*2048+   9, 
  25*2048+  42,   45*2048+  43,   45*2048+  44,   45*2048+  45,   12*2048+  46,   24*2048+  47,   40*2048+  48,   27*2048+  49,   45*2048+  50,   45*2048+  51, 
  45*2048+  99,   32*2048+ 100,   45*2048+ 101,   45*2048+ 102,   33*2048+ 103,   25*2048+ 104,   17*2048+ 105,   13*2048+ 106,   45*2048+ 107,   45*2048+ 108, 
  45*2048+ 132,   45*2048+ 133,   27*2048+ 134,   43*2048+ 135,   18*2048+ 136,   17*2048+ 137,   34*2048+ 138,   15*2048+ 139,   45*2048+ 140,   45*2048+ 141, 
  28*2048+ 174,   25*2048+ 175,   45*2048+ 176,   45*2048+ 177,   45*2048+ 178,   12*2048+ 179,   24*2048+ 180,   40*2048+ 181,   45*2048+ 182,   45*2048+ 183, 
  45*2048+ 231,   32*2048+ 232,   45*2048+ 233,   45*2048+ 234,   33*2048+ 235,   25*2048+ 236,   17*2048+ 237,   13*2048+ 238,   45*2048+ 239,   45*2048+ 240, 
  18*2048+ 264,   35*2048+ 265,   16*2048+ 266,   45*2048+ 267,   45*2048+ 268,   27*2048+ 269,   43*2048+ 270,   18*2048+ 271,   45*2048+ 272,   45*2048+ 273, 
  25*2048+ 306,   41*2048+ 307,   28*2048+ 308,   25*2048+ 309,   45*2048+ 310,   45*2048+ 311,   45*2048+ 312,   12*2048+ 313,   45*2048+ 314,   45*2048+ 315, 
  45*2048+ 363,   32*2048+ 364,   45*2048+ 365,   45*2048+ 366,   33*2048+ 367,   25*2048+ 368,   17*2048+ 369,   13*2048+ 370,   45*2048+ 371,   45*2048+ 372, 
  44*2048+ 396,   19*2048+ 397,   18*2048+ 398,   35*2048+ 399,   16*2048+ 400,   45*2048+ 401,   45*2048+ 402,   27*2048+ 403,   45*2048+ 404,   45*2048+ 405, 
  13*2048+ 438,   25*2048+ 439,   41*2048+ 440,   28*2048+ 441,   25*2048+ 442,   45*2048+ 443,   45*2048+ 444,   45*2048+ 445,   45*2048+ 446,   45*2048+ 447, 
  18*2048+ 495,   14*2048+ 496,   45*2048+ 497,   32*2048+ 498,   45*2048+ 499,   45*2048+ 500,   33*2048+ 501,   25*2048+ 502,   45*2048+ 503,   45*2048+ 504, 
  44*2048+ 528,   19*2048+ 529,   18*2048+ 530,   35*2048+ 531,   16*2048+ 532,   45*2048+ 533,   45*2048+ 534,   27*2048+ 535,   45*2048+ 536,   45*2048+ 537, 
  13*2048+ 570,   25*2048+ 571,   41*2048+ 572,   28*2048+ 573,   25*2048+ 574,   45*2048+ 575,   45*2048+ 576,   45*2048+ 577,   45*2048+ 578,   45*2048+ 579, 
  26*2048+ 627,   18*2048+ 628,   14*2048+ 629,   45*2048+ 630,   32*2048+ 631,   45*2048+ 632,   45*2048+ 633,   33*2048+ 634,   45*2048+ 635,   45*2048+ 636, 
  44*2048+ 660,   19*2048+ 661,   18*2048+ 662,   35*2048+ 663,   16*2048+ 664,   45*2048+ 665,   45*2048+ 666,   27*2048+ 667,   45*2048+ 668,   45*2048+ 669, 
  13*2048+ 702,   25*2048+ 703,   41*2048+ 704,   28*2048+ 705,   25*2048+ 706,   45*2048+ 707,   45*2048+ 708,   45*2048+ 709,   45*2048+ 710,   45*2048+ 711, 
  26*2048+ 759,   18*2048+ 760,   14*2048+ 761,   45*2048+ 762,   32*2048+ 763,   45*2048+ 764,   45*2048+ 765,   33*2048+ 766,   45*2048+ 767,   45*2048+ 768, 
  44*2048+ 792,   19*2048+ 793,   18*2048+ 794,   35*2048+ 795,   16*2048+ 796,   45*2048+ 797,   45*2048+ 798,   27*2048+ 799,   45*2048+ 800,   45*2048+ 801, 
  13*2048+ 834,   25*2048+ 835,   41*2048+ 836,   28*2048+ 837,   25*2048+ 838,   45*2048+ 839,   45*2048+ 840,   45*2048+ 841,   45*2048+ 842,   45*2048+ 843, 
  34*2048+ 891,   26*2048+ 892,   18*2048+ 893,   14*2048+ 894,   45*2048+ 895,   32*2048+ 896,   45*2048+ 897,   45*2048+ 898,   45*2048+ 899,   45*2048+ 900, 
  28*2048+ 924,   44*2048+ 925,   19*2048+ 926,   18*2048+ 927,   35*2048+ 928,   16*2048+ 929,   45*2048+ 930,   45*2048+ 931,   45*2048+ 932,   45*2048+ 933, 
  13*2048+ 966,   25*2048+ 967,   41*2048+ 968,   28*2048+ 969,   25*2048+ 970,   45*2048+ 971,   45*2048+ 972,   45*2048+ 973,   45*2048+ 974,   45*2048+ 975, 
  34*2048+1023,   26*2048+1024,   18*2048+1025,   14*2048+1026,   45*2048+1027,   32*2048+1028,   45*2048+1029,   45*2048+1030,   45*2048+1031,   45*2048+1032, 
  45*2048+  22,   45*2048+  23,    5*2048+  24,   39*2048+  25,   38*2048+  26,   39*2048+  27,   31*2048+  28,   34*2048+  29,   33*2048+  30,   45*2048+  31,   45*2048+  32, 
  45*2048+  65,   45*2048+  66,   45*2048+  67,   43*2048+  68,   16*2048+  69,   33*2048+  70,   11*2048+  71,   21*2048+  72,   29*2048+  73,   45*2048+  74,   45*2048+  75, 
  45*2048+  88,   45*2048+  89,   45*2048+  90,   31*2048+  91,    7*2048+  92,   19*2048+  93,    1*2048+  94,   23*2048+  95,   33*2048+  96,   45*2048+  97,   45*2048+  98, 
  45*2048+ 109,    4*2048+ 110,   45*2048+ 111,   45*2048+ 112,   40*2048+ 113,   27*2048+ 114,   26*2048+ 115,    6*2048+ 116,   43*2048+ 117,   45*2048+ 118,   45*2048+ 119, 
  34*2048+ 154,   45*2048+ 155,   45*2048+ 156,    5*2048+ 157,   39*2048+ 158,   38*2048+ 159,   39*2048+ 160,   31*2048+ 161,   34*2048+ 162,   45*2048+ 163,   45*2048+ 164, 
  30*2048+ 197,   45*2048+ 198,   45*2048+ 199,   45*2048+ 200,   43*2048+ 201,   16*2048+ 202,   33*2048+ 203,   11*2048+ 204,   21*2048+ 205,   45*2048+ 206,   45*2048+ 207, 
  45*2048+ 220,   45*2048+ 221,   45*2048+ 222,   31*2048+ 223,    7*2048+ 224,   19*2048+ 225,    1*2048+ 226,   23*2048+ 227,   33*2048+ 228,   45*2048+ 229,   45*2048+ 230, 
  45*2048+ 241,    4*2048+ 242,   45*2048+ 243,   45*2048+ 244,   40*2048+ 245,   27*2048+ 246,   26*2048+ 247,    6*2048+ 248,   43*2048+ 249,   45*2048+ 250,   45*2048+ 251, 
  35*2048+ 286,   34*2048+ 287,   45*2048+ 288,   45*2048+ 289,    5*2048+ 290,   39*2048+ 291,   38*2048+ 292,   39*2048+ 293,   31*2048+ 294,   45*2048+ 295,   45*2048+ 296, 
  12*2048+ 329,   22*2048+ 330,   30*2048+ 331,   45*2048+ 332,   45*2048+ 333,   45*2048+ 334,   43*2048+ 335,   16*2048+ 336,   33*2048+ 337,   45*2048+ 338,   45*2048+ 339, 
  34*2048+ 352,   45*2048+ 353,   45*2048+ 354,   45*2048+ 355,   31*2048+ 356,    7*2048+ 357,   19*2048+ 358,    1*2048+ 359,   23*2048+ 360,   45*2048+ 361,   45*2048+ 362, 
  45*2048+ 373,    4*2048+ 374,   45*2048+ 375,   45*2048+ 376,   40*2048+ 377,   27*2048+ 378,   26*2048+ 379,    6*2048+ 380,   43*2048+ 381,   45*2048+ 382,   45*2048+ 383, 
  35*2048+ 418,   34*2048+ 419,   45*2048+ 420,   45*2048+ 421,    5*2048+ 422,   39*2048+ 423,   38*2048+ 424,   39*2048+ 425,   31*2048+ 426,   45*2048+ 427,   45*2048+ 428, 
  12*2048+ 461,   22*2048+ 462,   30*2048+ 463,   45*2048+ 464,   45*2048+ 465,   45*2048+ 466,   43*2048+ 467,   16*2048+ 468,   33*2048+ 469,   45*2048+ 470,   45*2048+ 471, 
  24*2048+ 484,   34*2048+ 485,   45*2048+ 486,   45*2048+ 487,   45*2048+ 488,   31*2048+ 489,    7*2048+ 490,   19*2048+ 491,    1*2048+ 492,   45*2048+ 493,   45*2048+ 494, 
  27*2048+ 505,    7*2048+ 506,   44*2048+ 507,   45*2048+ 508,    4*2048+ 509,   45*2048+ 510,   45*2048+ 511,   40*2048+ 512,   27*2048+ 513,   45*2048+ 514,   45*2048+ 515, 
  32*2048+ 550,   35*2048+ 551,   34*2048+ 552,   45*2048+ 553,   45*2048+ 554,    5*2048+ 555,   39*2048+ 556,   38*2048+ 557,   39*2048+ 558,   45*2048+ 559,   45*2048+ 560, 
  17*2048+ 593,   34*2048+ 594,   12*2048+ 595,   22*2048+ 596,   30*2048+ 597,   45*2048+ 598,   45*2048+ 599,   45*2048+ 600,   43*2048+ 601,   45*2048+ 602,   45*2048+ 603, 
   2*2048+ 616,   24*2048+ 617,   34*2048+ 618,   45*2048+ 619,   45*2048+ 620,   45*2048+ 621,   31*2048+ 622,    7*2048+ 623,   19*2048+ 624,   45*2048+ 625,   45*2048+ 626, 
  28*2048+ 637,   27*2048+ 638,    7*2048+ 639,   44*2048+ 640,   45*2048+ 641,    4*2048+ 642,   45*2048+ 643,   45*2048+ 644,   40*2048+ 645,   45*2048+ 646,   45*2048+ 647, 
  39*2048+ 682,   40*2048+ 683,   32*2048+ 684,   35*2048+ 685,   34*2048+ 686,   45*2048+ 687,   45*2048+ 688,    5*2048+ 689,   39*2048+ 690,   45*2048+ 691,   45*2048+ 692, 
  17*2048+ 725,   34*2048+ 726,   12*2048+ 727,   22*2048+ 728,   30*2048+ 729,   45*2048+ 730,   45*2048+ 731,   45*2048+ 732,   43*2048+ 733,   45*2048+ 734,   45*2048+ 735, 
   2*2048+ 748,   24*2048+ 749,   34*2048+ 750,   45*2048+ 751,   45*2048+ 752,   45*2048+ 753,   31*2048+ 754,    7*2048+ 755,   19*2048+ 756,   45*2048+ 757,   45*2048+ 758, 
  28*2048+ 769,   27*2048+ 770,    7*2048+ 771,   44*2048+ 772,   45*2048+ 773,    4*2048+ 774,   45*2048+ 775,   45*2048+ 776,   40*2048+ 777,   45*2048+ 778,   45*2048+ 779, 
  40*2048+ 814,   39*2048+ 815,   40*2048+ 816,   32*2048+ 817,   35*2048+ 818,   34*2048+ 819,   45*2048+ 820,   45*2048+ 821,    5*2048+ 822,   45*2048+ 823,   45*2048+ 824, 
  44*2048+ 857,   17*2048+ 858,   34*2048+ 859,   12*2048+ 860,   22*2048+ 861,   30*2048+ 862,   45*2048+ 863,   45*2048+ 864,   45*2048+ 865,   45*2048+ 866,   45*2048+ 867, 
  32*2048+ 880,    8*2048+ 881,   20*2048+ 882,    2*2048+ 883,   24*2048+ 884,   34*2048+ 885,   45*2048+ 886,   45*2048+ 887,   45*2048+ 888,   45*2048+ 889,   45*2048+ 890, 
  28*2048+ 901,   27*2048+ 902,    7*2048+ 903,   44*2048+ 904,   45*2048+ 905,    4*2048+ 906,   45*2048+ 907,   45*2048+ 908,   40*2048+ 909,   45*2048+ 910,   45*2048+ 911, 
   6*2048+ 946,   40*2048+ 947,   39*2048+ 948,   40*2048+ 949,   32*2048+ 950,   35*2048+ 951,   34*2048+ 952,   45*2048+ 953,   45*2048+ 954,   45*2048+ 955,   45*2048+ 956, 
  44*2048+ 989,   17*2048+ 990,   34*2048+ 991,   12*2048+ 992,   22*2048+ 993,   30*2048+ 994,   45*2048+ 995,   45*2048+ 996,   45*2048+ 997,   45*2048+ 998,   45*2048+ 999, 
  32*2048+1012,    8*2048+1013,   20*2048+1014,    2*2048+1015,   24*2048+1016,   34*2048+1017,   45*2048+1018,   45*2048+1019,   45*2048+1020,   45*2048+1021,   45*2048+1022, 
  41*2048+1033,   28*2048+1034,   27*2048+1035,    7*2048+1036,   44*2048+1037,   45*2048+1038,    4*2048+1039,   45*2048+1040,   45*2048+1041,   45*2048+1042,   45*2048+1043, 
   2*2048+  10,   45*2048+  11,   45*2048+  12,   10*2048+  13,   26*2048+  14,   34*2048+  15,   34*2048+  16,   24*2048+  17,    9*2048+  18,    1*2048+  19,   45*2048+  20,   45*2048+  21, 
  45*2048+  76,   45*2048+  77,   13*2048+  78,   45*2048+  79,    3*2048+  80,    1*2048+  81,   13*2048+  82,   34*2048+  83,   21*2048+  84,   20*2048+  85,   45*2048+  86,   45*2048+  87, 
  38*2048+ 120,   45*2048+ 121,   45*2048+ 122,   45*2048+ 123,   25*2048+ 124,   30*2048+ 125,   12*2048+ 126,   34*2048+ 127,   30*2048+ 128,   22*2048+ 129,   45*2048+ 130,   45*2048+ 131, 
  10*2048+ 142,    2*2048+ 143,    2*2048+ 144,   45*2048+ 145,   45*2048+ 146,   10*2048+ 147,   26*2048+ 148,   34*2048+ 149,   34*2048+ 150,   24*2048+ 151,   45*2048+ 152,   45*2048+ 153, 
  21*2048+ 208,   45*2048+ 209,   45*2048+ 210,   13*2048+ 211,   45*2048+ 212,    3*2048+ 213,    1*2048+ 214,   13*2048+ 215,   34*2048+ 216,   21*2048+ 217,   45*2048+ 218,   45*2048+ 219, 
  23*2048+ 252,   38*2048+ 253,   45*2048+ 254,   45*2048+ 255,   45*2048+ 256,   25*2048+ 257,   30*2048+ 258,   12*2048+ 259,   34*2048+ 260,   30*2048+ 261,   45*2048+ 262,   45*2048+ 263, 
  25*2048+ 274,   10*2048+ 275,    2*2048+ 276,    2*2048+ 277,   45*2048+ 278,   45*2048+ 279,   10*2048+ 280,   26*2048+ 281,   34*2048+ 282,   34*2048+ 283,   45*2048+ 284,   45*2048+ 285, 
  22*2048+ 340,   21*2048+ 341,   45*2048+ 342,   45*2048+ 343,   13*2048+ 344,   45*2048+ 345,    3*2048+ 346,    1*2048+ 347,   13*2048+ 348,   34*2048+ 349,   45*2048+ 350,   45*2048+ 351, 
  13*2048+ 384,   35*2048+ 385,   31*2048+ 386,   23*2048+ 387,   38*2048+ 388,   45*2048+ 389,   45*2048+ 390,   45*2048+ 391,   25*2048+ 392,   30*2048+ 393,   45*2048+ 394,   45*2048+ 395, 
  35*2048+ 406,   25*2048+ 407,   10*2048+ 408,    2*2048+ 409,    2*2048+ 410,   45*2048+ 411,   45*2048+ 412,   10*2048+ 413,   26*2048+ 414,   34*2048+ 415,   45*2048+ 416,   45*2048+ 417, 
  22*2048+ 472,   21*2048+ 473,   45*2048+ 474,   45*2048+ 475,   13*2048+ 476,   45*2048+ 477,    3*2048+ 478,    1*2048+ 479,   13*2048+ 480,   34*2048+ 481,   45*2048+ 482,   45*2048+ 483, 
  13*2048+ 516,   35*2048+ 517,   31*2048+ 518,   23*2048+ 519,   38*2048+ 520,   45*2048+ 521,   45*2048+ 522,   45*2048+ 523,   25*2048+ 524,   30*2048+ 525,   45*2048+ 526,   45*2048+ 527, 
  35*2048+ 538,   35*2048+ 539,   25*2048+ 540,   10*2048+ 541,    2*2048+ 542,    2*2048+ 543,   45*2048+ 544,   45*2048+ 545,   10*2048+ 546,   26*2048+ 547,   45*2048+ 548,   45*2048+ 549, 
  14*2048+ 604,   35*2048+ 605,   22*2048+ 606,   21*2048+ 607,   45*2048+ 608,   45*2048+ 609,   13*2048+ 610,   45*2048+ 611,    3*2048+ 612,    1*2048+ 613,   45*2048+ 614,   45*2048+ 615, 
  13*2048+ 648,   35*2048+ 649,   31*2048+ 650,   23*2048+ 651,   38*2048+ 652,   45*2048+ 653,   45*2048+ 654,   45*2048+ 655,   25*2048+ 656,   30*2048+ 657,   45*2048+ 658,   45*2048+ 659, 
  35*2048+ 670,   35*2048+ 671,   25*2048+ 672,   10*2048+ 673,    2*2048+ 674,    2*2048+ 675,   45*2048+ 676,   45*2048+ 677,   10*2048+ 678,   26*2048+ 679,   45*2048+ 680,   45*2048+ 681, 
  14*2048+ 736,   35*2048+ 737,   22*2048+ 738,   21*2048+ 739,   45*2048+ 740,   45*2048+ 741,   13*2048+ 742,   45*2048+ 743,    3*2048+ 744,    1*2048+ 745,   45*2048+ 746,   45*2048+ 747, 
  31*2048+ 780,   13*2048+ 781,   35*2048+ 782,   31*2048+ 783,   23*2048+ 784,   38*2048+ 785,   45*2048+ 786,   45*2048+ 787,   45*2048+ 788,   25*2048+ 789,   45*2048+ 790,   45*2048+ 791, 
  27*2048+ 802,   35*2048+ 803,   35*2048+ 804,   25*2048+ 805,   10*2048+ 806,    2*2048+ 807,    2*2048+ 808,   45*2048+ 809,   45*2048+ 810,   10*2048+ 811,   45*2048+ 812,   45*2048+ 813, 
   2*2048+ 868,   14*2048+ 869,   35*2048+ 870,   22*2048+ 871,   21*2048+ 872,   45*2048+ 873,   45*2048+ 874,   13*2048+ 875,   45*2048+ 876,    3*2048+ 877,   45*2048+ 878,   45*2048+ 879, 
  26*2048+ 912,   31*2048+ 913,   13*2048+ 914,   35*2048+ 915,   31*2048+ 916,   23*2048+ 917,   38*2048+ 918,   45*2048+ 919,   45*2048+ 920,   45*2048+ 921,   45*2048+ 922,   45*2048+ 923, 
  27*2048+ 934,   35*2048+ 935,   35*2048+ 936,   25*2048+ 937,   10*2048+ 938,    2*2048+ 939,    2*2048+ 940,   45*2048+ 941,   45*2048+ 942,   10*2048+ 943,   45*2048+ 944,   45*2048+ 945, 
   4*2048+1000,    2*2048+1001,   14*2048+1002,   35*2048+1003,   22*2048+1004,   21*2048+1005,   45*2048+1006,   45*2048+1007,   13*2048+1008,   45*2048+1009,   45*2048+1010,   45*2048+1011, 
  26*2048+1044,   31*2048+1045,   13*2048+1046,   35*2048+1047,   31*2048+1048,   23*2048+1049,   38*2048+1050,   45*2048+1051,   45*2048+1052,   45*2048+1053,   45*2048+1054,   45*2048+1055, 
  45*2048+  52,   45*2048+  53,   45*2048+  54,   20*2048+  55,   17*2048+  56,    9*2048+  57,   26*2048+  58,    9*2048+  59,    6*2048+  60,   29*2048+  61,   37*2048+  62,   45*2048+  63,   45*2048+  64, 
  45*2048+ 184,   45*2048+ 185,   45*2048+ 186,   20*2048+ 187,   17*2048+ 188,    9*2048+ 189,   26*2048+ 190,    9*2048+ 191,    6*2048+ 192,   29*2048+ 193,   37*2048+ 194,   45*2048+ 195,   45*2048+ 196, 
  45*2048+ 316,   45*2048+ 317,   45*2048+ 318,   20*2048+ 319,   17*2048+ 320,    9*2048+ 321,   26*2048+ 322,    9*2048+ 323,    6*2048+ 324,   29*2048+ 325,   37*2048+ 326,   45*2048+ 327,   45*2048+ 328, 
  30*2048+ 448,   38*2048+ 449,   45*2048+ 450,   45*2048+ 451,   45*2048+ 452,   20*2048+ 453,   17*2048+ 454,    9*2048+ 455,   26*2048+ 456,    9*2048+ 457,    6*2048+ 458,   45*2048+ 459,   45*2048+ 460, 
  30*2048+ 580,   38*2048+ 581,   45*2048+ 582,   45*2048+ 583,   45*2048+ 584,   20*2048+ 585,   17*2048+ 586,    9*2048+ 587,   26*2048+ 588,    9*2048+ 589,    6*2048+ 590,   45*2048+ 591,   45*2048+ 592, 
  30*2048+ 712,   38*2048+ 713,   45*2048+ 714,   45*2048+ 715,   45*2048+ 716,   20*2048+ 717,   17*2048+ 718,    9*2048+ 719,   26*2048+ 720,    9*2048+ 721,    6*2048+ 722,   45*2048+ 723,   45*2048+ 724, 
  10*2048+ 844,    7*2048+ 845,   30*2048+ 846,   38*2048+ 847,   45*2048+ 848,   45*2048+ 849,   45*2048+ 850,   20*2048+ 851,   17*2048+ 852,    9*2048+ 853,   26*2048+ 854,   45*2048+ 855,   45*2048+ 856, 
  18*2048+ 976,   10*2048+ 977,   27*2048+ 978,   10*2048+ 979,    7*2048+ 980,   30*2048+ 981,   38*2048+ 982,   45*2048+ 983,   45*2048+ 984,   45*2048+ 985,   20*2048+ 986,   45*2048+ 987,   45*2048+ 988, 

  45*2048+  12,   45*2048+  13,   45*2048+  14,   33*2048+  15,   27*2048+  16,   11*2048+  17,   43*2048+  18,   21*2048+  19,   40*2048+  20,   45*2048+  21,   45*2048+  22, 
  41*2048+ 137,   45*2048+ 138,   45*2048+ 139,   45*2048+ 140,   33*2048+ 141,   27*2048+ 142,   11*2048+ 143,   43*2048+ 144,   21*2048+ 145,   45*2048+ 146,   45*2048+ 147, 
  41*2048+ 262,   45*2048+ 263,   45*2048+ 264,   45*2048+ 265,   33*2048+ 266,   27*2048+ 267,   11*2048+ 268,   43*2048+ 269,   21*2048+ 270,   45*2048+ 271,   45*2048+ 272, 
  41*2048+ 387,   45*2048+ 388,   45*2048+ 389,   45*2048+ 390,   33*2048+ 391,   27*2048+ 392,   11*2048+ 393,   43*2048+ 394,   21*2048+ 395,   45*2048+ 396,   45*2048+ 397, 
  44*2048+ 512,   22*2048+ 513,   41*2048+ 514,   45*2048+ 515,   45*2048+ 516,   45*2048+ 517,   33*2048+ 518,   27*2048+ 519,   11*2048+ 520,   45*2048+ 521,   45*2048+ 522, 
  44*2048+ 637,   22*2048+ 638,   41*2048+ 639,   45*2048+ 640,   45*2048+ 641,   45*2048+ 642,   33*2048+ 643,   27*2048+ 644,   11*2048+ 645,   45*2048+ 646,   45*2048+ 647, 
  28*2048+ 762,   12*2048+ 763,   44*2048+ 764,   22*2048+ 765,   41*2048+ 766,   45*2048+ 767,   45*2048+ 768,   45*2048+ 769,   33*2048+ 770,   45*2048+ 771,   45*2048+ 772, 
  34*2048+ 887,   28*2048+ 888,   12*2048+ 889,   44*2048+ 890,   22*2048+ 891,   41*2048+ 892,   45*2048+ 893,   45*2048+ 894,   45*2048+ 895,   45*2048+ 896,   45*2048+ 897, 
  45*2048+   0,   45*2048+   1,    4*2048+   2,   45*2048+   3,   42*2048+   4,   22*2048+   5,   18*2048+   6,    1*2048+   7,    4*2048+   8,   24*2048+   9,   45*2048+  10,   44*2048+  11, 
  45*2048+  36,   45*2048+  37,   45*2048+  38,    4*2048+  39,   42*2048+  40,   41*2048+  41,   11*2048+  42,   27*2048+  43,   40*2048+  44,   13*2048+  45,   45*2048+  46,   45*2048+  47, 
  45*2048+  48,   45*2048+  49,   45*2048+  50,   10*2048+  51,   25*2048+  52,   10*2048+  53,   19*2048+  54,    6*2048+  55,   42*2048+  56,   43*2048+  57,   45*2048+  58,   45*2048+  59, 
   5*2048+ 125,   25*2048+ 126,   45*2048+ 127,   45*2048+ 128,    4*2048+ 129,   45*2048+ 130,   42*2048+ 131,   22*2048+ 132,   18*2048+ 133,    1*2048+ 134,   45*2048+ 135,   45*2048+ 136, 
  14*2048+ 161,   45*2048+ 162,   45*2048+ 163,   45*2048+ 164,    4*2048+ 165,   42*2048+ 166,   41*2048+ 167,   11*2048+ 168,   27*2048+ 169,   40*2048+ 170,   45*2048+ 171,   45*2048+ 172, 
  44*2048+ 173,   45*2048+ 174,   45*2048+ 175,   45*2048+ 176,   10*2048+ 177,   25*2048+ 178,   10*2048+ 179,   19*2048+ 180,    6*2048+ 181,   42*2048+ 182,   45*2048+ 183,   45*2048+ 184, 
   2*2048+ 250,    5*2048+ 251,   25*2048+ 252,   45*2048+ 253,   45*2048+ 254,    4*2048+ 255,   45*2048+ 256,   42*2048+ 257,   22*2048+ 258,   18*2048+ 259,   45*2048+ 260,   45*2048+ 261, 
  12*2048+ 286,   28*2048+ 287,   41*2048+ 288,   14*2048+ 289,   45*2048+ 290,   45*2048+ 291,   45*2048+ 292,    4*2048+ 293,   42*2048+ 294,   41*2048+ 295,   45*2048+ 296,   45*2048+ 297, 
  43*2048+ 298,   44*2048+ 299,   45*2048+ 300,   45*2048+ 301,   45*2048+ 302,   10*2048+ 303,   25*2048+ 304,   10*2048+ 305,   19*2048+ 306,    6*2048+ 307,   45*2048+ 308,   45*2048+ 309, 
  19*2048+ 375,    2*2048+ 376,    5*2048+ 377,   25*2048+ 378,   45*2048+ 379,   45*2048+ 380,    4*2048+ 381,   45*2048+ 382,   42*2048+ 383,   22*2048+ 384,   45*2048+ 385,   45*2048+ 386, 
  12*2048+ 411,   28*2048+ 412,   41*2048+ 413,   14*2048+ 414,   45*2048+ 415,   45*2048+ 416,   45*2048+ 417,    4*2048+ 418,   42*2048+ 419,   41*2048+ 420,   45*2048+ 421,   45*2048+ 422, 
  20*2048+ 423,    7*2048+ 424,   43*2048+ 425,   44*2048+ 426,   45*2048+ 427,   45*2048+ 428,   45*2048+ 429,   10*2048+ 430,   25*2048+ 431,   10*2048+ 432,   45*2048+ 433,   45*2048+ 434, 
  23*2048+ 500,   19*2048+ 501,    2*2048+ 502,    5*2048+ 503,   25*2048+ 504,   45*2048+ 505,   45*2048+ 506,    4*2048+ 507,   45*2048+ 508,   42*2048+ 509,   45*2048+ 510,   45*2048+ 511, 
  42*2048+ 536,   12*2048+ 537,   28*2048+ 538,   41*2048+ 539,   14*2048+ 540,   45*2048+ 541,   45*2048+ 542,   45*2048+ 543,    4*2048+ 544,   42*2048+ 545,   45*2048+ 546,   45*2048+ 547, 
  20*2048+ 548,    7*2048+ 549,   43*2048+ 550,   44*2048+ 551,   45*2048+ 552,   45*2048+ 553,   45*2048+ 554,   10*2048+ 555,   25*2048+ 556,   10*2048+ 557,   45*2048+ 558,   45*2048+ 559, 
  23*2048+ 625,   19*2048+ 626,    2*2048+ 627,    5*2048+ 628,   25*2048+ 629,   45*2048+ 630,   45*2048+ 631,    4*2048+ 632,   45*2048+ 633,   42*2048+ 634,   45*2048+ 635,   45*2048+ 636, 
  42*2048+ 661,   12*2048+ 662,   28*2048+ 663,   41*2048+ 664,   14*2048+ 665,   45*2048+ 666,   45*2048+ 667,   45*2048+ 668,    4*2048+ 669,   42*2048+ 670,   45*2048+ 671,   45*2048+ 672, 
  11*2048+ 673,   20*2048+ 674,    7*2048+ 675,   43*2048+ 676,   44*2048+ 677,   45*2048+ 678,   45*2048+ 679,   45*2048+ 680,   10*2048+ 681,   25*2048+ 682,   45*2048+ 683,   45*2048+ 684, 
  23*2048+ 750,   19*2048+ 751,    2*2048+ 752,    5*2048+ 753,   25*2048+ 754,   45*2048+ 755,   45*2048+ 756,    4*2048+ 757,   45*2048+ 758,   42*2048+ 759,   45*2048+ 760,   45*2048+ 761, 
  42*2048+ 786,   12*2048+ 787,   28*2048+ 788,   41*2048+ 789,   14*2048+ 790,   45*2048+ 791,   45*2048+ 792,   45*2048+ 793,    4*2048+ 794,   42*2048+ 795,   45*2048+ 796,   45*2048+ 797, 
  26*2048+ 798,   11*2048+ 799,   20*2048+ 800,    7*2048+ 801,   43*2048+ 802,   44*2048+ 803,   45*2048+ 804,   45*2048+ 805,   45*2048+ 806,   10*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  43*2048+ 875,   23*2048+ 876,   19*2048+ 877,    2*2048+ 878,    5*2048+ 879,   25*2048+ 880,   45*2048+ 881,   45*2048+ 882,    4*2048+ 883,   45*2048+ 884,   45*2048+ 885,   45*2048+ 886, 
  42*2048+ 911,   12*2048+ 912,   28*2048+ 913,   41*2048+ 914,   14*2048+ 915,   45*2048+ 916,   45*2048+ 917,   45*2048+ 918,    4*2048+ 919,   42*2048+ 920,   45*2048+ 921,   45*2048+ 922, 
  11*2048+ 923,   26*2048+ 924,   11*2048+ 925,   20*2048+ 926,    7*2048+ 927,   43*2048+ 928,   44*2048+ 929,   45*2048+ 930,   45*2048+ 931,   45*2048+ 932,   45*2048+ 933,   45*2048+ 934, 
  45*2048+  23,   45*2048+  24,   36*2048+  25,   45*2048+  26,   13*2048+  27,   34*2048+  28,   42*2048+  29,   37*2048+  30,   23*2048+  31,   16*2048+  32,    0*2048+  33,   45*2048+  34,   45*2048+  35, 
  45*2048+  60,   45*2048+  61,   45*2048+  62,   45*2048+  63,   39*2048+  64,   33*2048+  65,   11*2048+  66,   25*2048+  67,   19*2048+  68,    0*2048+  69,   21*2048+  70,   45*2048+  71,   45*2048+  72, 
  45*2048+  73,   45*2048+  74,   45*2048+  75,   45*2048+  76,   38*2048+  77,   42*2048+  78,   23*2048+  79,   40*2048+  80,   16*2048+  81,   18*2048+  82,   33*2048+  83,   45*2048+  84,   45*2048+  85, 
  45*2048+  86,   36*2048+  87,   45*2048+  88,   45*2048+  89,   45*2048+  90,   30*2048+  91,   41*2048+  92,   27*2048+  93,   26*2048+  94,   10*2048+  95,   20*2048+  96,   45*2048+  97,   45*2048+  98, 
  45*2048+  99,   45*2048+ 100,   45*2048+ 101,   43*2048+ 102,   45*2048+ 103,   32*2048+ 104,    2*2048+ 105,   19*2048+ 106,    6*2048+ 107,   16*2048+ 108,   30*2048+ 109,   45*2048+ 110,   45*2048+ 111, 
  45*2048+ 112,    9*2048+ 113,   45*2048+ 114,   45*2048+ 115,   45*2048+ 116,    7*2048+ 117,   14*2048+ 118,   28*2048+ 119,   12*2048+ 120,   31*2048+ 121,   19*2048+ 122,   45*2048+ 123,   45*2048+ 124, 
  45*2048+ 148,   45*2048+ 149,   36*2048+ 150,   45*2048+ 151,   13*2048+ 152,   34*2048+ 153,   42*2048+ 154,   37*2048+ 155,   23*2048+ 156,   16*2048+ 157,    0*2048+ 158,   45*2048+ 159,   45*2048+ 160, 
  22*2048+ 185,   45*2048+ 186,   45*2048+ 187,   45*2048+ 188,   45*2048+ 189,   39*2048+ 190,   33*2048+ 191,   11*2048+ 192,   25*2048+ 193,   19*2048+ 194,    0*2048+ 195,   45*2048+ 196,   45*2048+ 197, 
  34*2048+ 198,   45*2048+ 199,   45*2048+ 200,   45*2048+ 201,   45*2048+ 202,   38*2048+ 203,   42*2048+ 204,   23*2048+ 205,   40*2048+ 206,   16*2048+ 207,   18*2048+ 208,   45*2048+ 209,   45*2048+ 210, 
  45*2048+ 211,   36*2048+ 212,   45*2048+ 213,   45*2048+ 214,   45*2048+ 215,   30*2048+ 216,   41*2048+ 217,   27*2048+ 218,   26*2048+ 219,   10*2048+ 220,   20*2048+ 221,   45*2048+ 222,   45*2048+ 223, 
  45*2048+ 224,   45*2048+ 225,   45*2048+ 226,   43*2048+ 227,   45*2048+ 228,   32*2048+ 229,    2*2048+ 230,   19*2048+ 231,    6*2048+ 232,   16*2048+ 233,   30*2048+ 234,   45*2048+ 235,   45*2048+ 236, 
  45*2048+ 237,    9*2048+ 238,   45*2048+ 239,   45*2048+ 240,   45*2048+ 241,    7*2048+ 242,   14*2048+ 243,   28*2048+ 244,   12*2048+ 245,   31*2048+ 246,   19*2048+ 247,   45*2048+ 248,   45*2048+ 249, 
   1*2048+ 273,   45*2048+ 274,   45*2048+ 275,   36*2048+ 276,   45*2048+ 277,   13*2048+ 278,   34*2048+ 279,   42*2048+ 280,   37*2048+ 281,   23*2048+ 282,   16*2048+ 283,   45*2048+ 284,   45*2048+ 285, 
  20*2048+ 310,    1*2048+ 311,   22*2048+ 312,   45*2048+ 313,   45*2048+ 314,   45*2048+ 315,   45*2048+ 316,   39*2048+ 317,   33*2048+ 318,   11*2048+ 319,   25*2048+ 320,   45*2048+ 321,   45*2048+ 322, 
  34*2048+ 323,   45*2048+ 324,   45*2048+ 325,   45*2048+ 326,   45*2048+ 327,   38*2048+ 328,   42*2048+ 329,   23*2048+ 330,   40*2048+ 331,   16*2048+ 332,   18*2048+ 333,   45*2048+ 334,   45*2048+ 335, 
  21*2048+ 336,   45*2048+ 337,   36*2048+ 338,   45*2048+ 339,   45*2048+ 340,   45*2048+ 341,   30*2048+ 342,   41*2048+ 343,   27*2048+ 344,   26*2048+ 345,   10*2048+ 346,   45*2048+ 347,   45*2048+ 348, 
  45*2048+ 349,   45*2048+ 350,   45*2048+ 351,   43*2048+ 352,   45*2048+ 353,   32*2048+ 354,    2*2048+ 355,   19*2048+ 356,    6*2048+ 357,   16*2048+ 358,   30*2048+ 359,   45*2048+ 360,   45*2048+ 361, 
  45*2048+ 362,    9*2048+ 363,   45*2048+ 364,   45*2048+ 365,   45*2048+ 366,    7*2048+ 367,   14*2048+ 368,   28*2048+ 369,   12*2048+ 370,   31*2048+ 371,   19*2048+ 372,   45*2048+ 373,   45*2048+ 374, 
  17*2048+ 398,    1*2048+ 399,   45*2048+ 400,   45*2048+ 401,   36*2048+ 402,   45*2048+ 403,   13*2048+ 404,   34*2048+ 405,   42*2048+ 406,   37*2048+ 407,   23*2048+ 408,   45*2048+ 409,   45*2048+ 410, 
  20*2048+ 435,    1*2048+ 436,   22*2048+ 437,   45*2048+ 438,   45*2048+ 439,   45*2048+ 440,   45*2048+ 441,   39*2048+ 442,   33*2048+ 443,   11*2048+ 444,   25*2048+ 445,   45*2048+ 446,   45*2048+ 447, 
  19*2048+ 448,   34*2048+ 449,   45*2048+ 450,   45*2048+ 451,   45*2048+ 452,   45*2048+ 453,   38*2048+ 454,   42*2048+ 455,   23*2048+ 456,   40*2048+ 457,   16*2048+ 458,   45*2048+ 459,   45*2048+ 460, 
  21*2048+ 461,   45*2048+ 462,   36*2048+ 463,   45*2048+ 464,   45*2048+ 465,   45*2048+ 466,   30*2048+ 467,   41*2048+ 468,   27*2048+ 469,   26*2048+ 470,   10*2048+ 471,   45*2048+ 472,   45*2048+ 473, 
  45*2048+ 474,   45*2048+ 475,   45*2048+ 476,   43*2048+ 477,   45*2048+ 478,   32*2048+ 479,    2*2048+ 480,   19*2048+ 481,    6*2048+ 482,   16*2048+ 483,   30*2048+ 484,   45*2048+ 485,   45*2048+ 486, 
  45*2048+ 487,    9*2048+ 488,   45*2048+ 489,   45*2048+ 490,   45*2048+ 491,    7*2048+ 492,   14*2048+ 493,   28*2048+ 494,   12*2048+ 495,   31*2048+ 496,   19*2048+ 497,   45*2048+ 498,   45*2048+ 499, 
  17*2048+ 523,    1*2048+ 524,   45*2048+ 525,   45*2048+ 526,   36*2048+ 527,   45*2048+ 528,   13*2048+ 529,   34*2048+ 530,   42*2048+ 531,   37*2048+ 532,   23*2048+ 533,   45*2048+ 534,   45*2048+ 535, 
  26*2048+ 560,   20*2048+ 561,    1*2048+ 562,   22*2048+ 563,   45*2048+ 564,   45*2048+ 565,   45*2048+ 566,   45*2048+ 567,   39*2048+ 568,   33*2048+ 569,   11*2048+ 570,   45*2048+ 571,   45*2048+ 572, 
  17*2048+ 573,   19*2048+ 574,   34*2048+ 575,   45*2048+ 576,   45*2048+ 577,   45*2048+ 578,   45*2048+ 579,   38*2048+ 580,   42*2048+ 581,   23*2048+ 582,   40*2048+ 583,   45*2048+ 584,   45*2048+ 585, 
  11*2048+ 586,   21*2048+ 587,   45*2048+ 588,   36*2048+ 589,   45*2048+ 590,   45*2048+ 591,   45*2048+ 592,   30*2048+ 593,   41*2048+ 594,   27*2048+ 595,   26*2048+ 596,   45*2048+ 597,   45*2048+ 598, 
  31*2048+ 599,   45*2048+ 600,   45*2048+ 601,   45*2048+ 602,   43*2048+ 603,   45*2048+ 604,   32*2048+ 605,    2*2048+ 606,   19*2048+ 607,    6*2048+ 608,   16*2048+ 609,   45*2048+ 610,   45*2048+ 611, 
  20*2048+ 612,   45*2048+ 613,    9*2048+ 614,   45*2048+ 615,   45*2048+ 616,   45*2048+ 617,    7*2048+ 618,   14*2048+ 619,   28*2048+ 620,   12*2048+ 621,   31*2048+ 622,   45*2048+ 623,   45*2048+ 624, 
  43*2048+ 648,   38*2048+ 649,   24*2048+ 650,   17*2048+ 651,    1*2048+ 652,   45*2048+ 653,   45*2048+ 654,   36*2048+ 655,   45*2048+ 656,   13*2048+ 657,   34*2048+ 658,   45*2048+ 659,   45*2048+ 660, 
  12*2048+ 685,   26*2048+ 686,   20*2048+ 687,    1*2048+ 688,   22*2048+ 689,   45*2048+ 690,   45*2048+ 691,   45*2048+ 692,   45*2048+ 693,   39*2048+ 694,   33*2048+ 695,   45*2048+ 696,   45*2048+ 697, 
  41*2048+ 698,   17*2048+ 699,   19*2048+ 700,   34*2048+ 701,   45*2048+ 702,   45*2048+ 703,   45*2048+ 704,   45*2048+ 705,   38*2048+ 706,   42*2048+ 707,   23*2048+ 708,   45*2048+ 709,   45*2048+ 710, 
  27*2048+ 711,   11*2048+ 712,   21*2048+ 713,   45*2048+ 714,   36*2048+ 715,   45*2048+ 716,   45*2048+ 717,   45*2048+ 718,   30*2048+ 719,   41*2048+ 720,   27*2048+ 721,   45*2048+ 722,   45*2048+ 723, 
  31*2048+ 724,   45*2048+ 725,   45*2048+ 726,   45*2048+ 727,   43*2048+ 728,   45*2048+ 729,   32*2048+ 730,    2*2048+ 731,   19*2048+ 732,    6*2048+ 733,   16*2048+ 734,   45*2048+ 735,   45*2048+ 736, 
  29*2048+ 737,   13*2048+ 738,   32*2048+ 739,   20*2048+ 740,   45*2048+ 741,    9*2048+ 742,   45*2048+ 743,   45*2048+ 744,   45*2048+ 745,    7*2048+ 746,   14*2048+ 747,   45*2048+ 748,   45*2048+ 749, 
  35*2048+ 773,   43*2048+ 774,   38*2048+ 775,   24*2048+ 776,   17*2048+ 777,    1*2048+ 778,   45*2048+ 779,   45*2048+ 780,   36*2048+ 781,   45*2048+ 782,   13*2048+ 783,   45*2048+ 784,   45*2048+ 785, 
  40*2048+ 810,   34*2048+ 811,   12*2048+ 812,   26*2048+ 813,   20*2048+ 814,    1*2048+ 815,   22*2048+ 816,   45*2048+ 817,   45*2048+ 818,   45*2048+ 819,   45*2048+ 820,   45*2048+ 821,   45*2048+ 822, 
  24*2048+ 823,   41*2048+ 824,   17*2048+ 825,   19*2048+ 826,   34*2048+ 827,   45*2048+ 828,   45*2048+ 829,   45*2048+ 830,   45*2048+ 831,   38*2048+ 832,   42*2048+ 833,   45*2048+ 834,   45*2048+ 835, 
  42*2048+ 836,   28*2048+ 837,   27*2048+ 838,   11*2048+ 839,   21*2048+ 840,   45*2048+ 841,   36*2048+ 842,   45*2048+ 843,   45*2048+ 844,   45*2048+ 845,   30*2048+ 846,   45*2048+ 847,   45*2048+ 848, 
   3*2048+ 849,   20*2048+ 850,    7*2048+ 851,   17*2048+ 852,   31*2048+ 853,   45*2048+ 854,   45*2048+ 855,   45*2048+ 856,   43*2048+ 857,   45*2048+ 858,   32*2048+ 859,   45*2048+ 860,   45*2048+ 861, 
  29*2048+ 862,   13*2048+ 863,   32*2048+ 864,   20*2048+ 865,   45*2048+ 866,    9*2048+ 867,   45*2048+ 868,   45*2048+ 869,   45*2048+ 870,    7*2048+ 871,   14*2048+ 872,   45*2048+ 873,   45*2048+ 874, 
  14*2048+ 898,   35*2048+ 899,   43*2048+ 900,   38*2048+ 901,   24*2048+ 902,   17*2048+ 903,    1*2048+ 904,   45*2048+ 905,   45*2048+ 906,   36*2048+ 907,   45*2048+ 908,   45*2048+ 909,   45*2048+ 910, 
  40*2048+ 935,   34*2048+ 936,   12*2048+ 937,   26*2048+ 938,   20*2048+ 939,    1*2048+ 940,   22*2048+ 941,   45*2048+ 942,   45*2048+ 943,   45*2048+ 944,   45*2048+ 945,   45*2048+ 946,   45*2048+ 947, 
  43*2048+ 948,   24*2048+ 949,   41*2048+ 950,   17*2048+ 951,   19*2048+ 952,   34*2048+ 953,   45*2048+ 954,   45*2048+ 955,   45*2048+ 956,   45*2048+ 957,   38*2048+ 958,   45*2048+ 959,   45*2048+ 960, 
  31*2048+ 961,   42*2048+ 962,   28*2048+ 963,   27*2048+ 964,   11*2048+ 965,   21*2048+ 966,   45*2048+ 967,   36*2048+ 968,   45*2048+ 969,   45*2048+ 970,   45*2048+ 971,   45*2048+ 972,   45*2048+ 973, 
  33*2048+ 974,    3*2048+ 975,   20*2048+ 976,    7*2048+ 977,   17*2048+ 978,   31*2048+ 979,   45*2048+ 980,   45*2048+ 981,   45*2048+ 982,   43*2048+ 983,   45*2048+ 984,   45*2048+ 985,   45*2048+ 986, 
   8*2048+ 987,   15*2048+ 988,   29*2048+ 989,   13*2048+ 990,   32*2048+ 991,   20*2048+ 992,   45*2048+ 993,    9*2048+ 994,   45*2048+ 995,   45*2048+ 996,   45*2048+ 997,   45*2048+ 998,   45*2048+ 999, 

  45*2048+   0,   12*2048+   1,   45*2048+   2,   45*2048+   3,   41*2048+   4,   45*2048+   5,   25*2048+   6,   18*2048+   7,   18*2048+   8,    9*2048+   9,    7*2048+  10,   27*2048+  11,    8*2048+  12,   25*2048+  13,   45*2048+  14,   44*2048+  15, 
  45*2048+  16,   45*2048+  17,   45*2048+  18,    8*2048+  19,   45*2048+  20,   44*2048+  21,   37*2048+  22,    7*2048+  23,   42*2048+  24,   25*2048+  25,   36*2048+  26,   43*2048+  27,   21*2048+  28,   25*2048+  29,   45*2048+  30,   45*2048+  31, 
  12*2048+  32,   45*2048+  33,   45*2048+  34,   45*2048+  35,   45*2048+  36,   15*2048+  37,   19*2048+  38,   43*2048+  39,    6*2048+  40,   22*2048+  41,   28*2048+  42,    9*2048+  43,   31*2048+  44,   17*2048+  45,   45*2048+  46,   45*2048+  47, 
  45*2048+  48,   45*2048+  49,   10*2048+  50,   45*2048+  51,   45*2048+  52,   45*2048+  53,   37*2048+  54,   32*2048+  55,    3*2048+  56,   38*2048+  57,   20*2048+  58,   37*2048+  59,   42*2048+  60,   43*2048+  61,   45*2048+  62,   45*2048+  63, 
  26*2048+ 137,   45*2048+ 138,   12*2048+ 139,   45*2048+ 140,   45*2048+ 141,   41*2048+ 142,   45*2048+ 143,   25*2048+ 144,   18*2048+ 145,   18*2048+ 146,    9*2048+ 147,    7*2048+ 148,   27*2048+ 149,    8*2048+ 150,   45*2048+ 151,   45*2048+ 152, 
  22*2048+ 153,   26*2048+ 154,   45*2048+ 155,   45*2048+ 156,   45*2048+ 157,    8*2048+ 158,   45*2048+ 159,   44*2048+ 160,   37*2048+ 161,    7*2048+ 162,   42*2048+ 163,   25*2048+ 164,   36*2048+ 165,   43*2048+ 166,   45*2048+ 167,   45*2048+ 168, 
  32*2048+ 169,   18*2048+ 170,   12*2048+ 171,   45*2048+ 172,   45*2048+ 173,   45*2048+ 174,   45*2048+ 175,   15*2048+ 176,   19*2048+ 177,   43*2048+ 178,    6*2048+ 179,   22*2048+ 180,   28*2048+ 181,    9*2048+ 182,   45*2048+ 183,   45*2048+ 184, 
  45*2048+ 185,   45*2048+ 186,   10*2048+ 187,   45*2048+ 188,   45*2048+ 189,   45*2048+ 190,   37*2048+ 191,   32*2048+ 192,    3*2048+ 193,   38*2048+ 194,   20*2048+ 195,   37*2048+ 196,   42*2048+ 197,   43*2048+ 198,   45*2048+ 199,   45*2048+ 200, 
  28*2048+ 274,    9*2048+ 275,   26*2048+ 276,   45*2048+ 277,   12*2048+ 278,   45*2048+ 279,   45*2048+ 280,   41*2048+ 281,   45*2048+ 282,   25*2048+ 283,   18*2048+ 284,   18*2048+ 285,    9*2048+ 286,    7*2048+ 287,   45*2048+ 288,   45*2048+ 289, 
  44*2048+ 290,   22*2048+ 291,   26*2048+ 292,   45*2048+ 293,   45*2048+ 294,   45*2048+ 295,    8*2048+ 296,   45*2048+ 297,   44*2048+ 298,   37*2048+ 299,    7*2048+ 300,   42*2048+ 301,   25*2048+ 302,   36*2048+ 303,   45*2048+ 304,   45*2048+ 305, 
  10*2048+ 306,   32*2048+ 307,   18*2048+ 308,   12*2048+ 309,   45*2048+ 310,   45*2048+ 311,   45*2048+ 312,   45*2048+ 313,   15*2048+ 314,   19*2048+ 315,   43*2048+ 316,    6*2048+ 317,   22*2048+ 318,   28*2048+ 319,   45*2048+ 320,   45*2048+ 321, 
  45*2048+ 322,   45*2048+ 323,   10*2048+ 324,   45*2048+ 325,   45*2048+ 326,   45*2048+ 327,   37*2048+ 328,   32*2048+ 329,    3*2048+ 330,   38*2048+ 331,   20*2048+ 332,   37*2048+ 333,   42*2048+ 334,   43*2048+ 335,   45*2048+ 336,   45*2048+ 337, 
  10*2048+ 411,    8*2048+ 412,   28*2048+ 413,    9*2048+ 414,   26*2048+ 415,   45*2048+ 416,   12*2048+ 417,   45*2048+ 418,   45*2048+ 419,   41*2048+ 420,   45*2048+ 421,   25*2048+ 422,   18*2048+ 423,   18*2048+ 424,   45*2048+ 425,   45*2048+ 426, 
  44*2048+ 427,   22*2048+ 428,   26*2048+ 429,   45*2048+ 430,   45*2048+ 431,   45*2048+ 432,    8*2048+ 433,   45*2048+ 434,   44*2048+ 435,   37*2048+ 436,    7*2048+ 437,   42*2048+ 438,   25*2048+ 439,   36*2048+ 440,   45*2048+ 441,   45*2048+ 442, 
  29*2048+ 443,   10*2048+ 444,   32*2048+ 445,   18*2048+ 446,   12*2048+ 447,   45*2048+ 448,   45*2048+ 449,   45*2048+ 450,   45*2048+ 451,   15*2048+ 452,   19*2048+ 453,   43*2048+ 454,    6*2048+ 455,   22*2048+ 456,   45*2048+ 457,   45*2048+ 458, 
  44*2048+ 459,   45*2048+ 460,   45*2048+ 461,   10*2048+ 462,   45*2048+ 463,   45*2048+ 464,   45*2048+ 465,   37*2048+ 466,   32*2048+ 467,    3*2048+ 468,   38*2048+ 469,   20*2048+ 470,   37*2048+ 471,   42*2048+ 472,   45*2048+ 473,   45*2048+ 474, 
  19*2048+ 548,   10*2048+ 549,    8*2048+ 550,   28*2048+ 551,    9*2048+ 552,   26*2048+ 553,   45*2048+ 554,   12*2048+ 555,   45*2048+ 556,   45*2048+ 557,   41*2048+ 558,   45*2048+ 559,   25*2048+ 560,   18*2048+ 561,   45*2048+ 562,   45*2048+ 563, 
  37*2048+ 564,   44*2048+ 565,   22*2048+ 566,   26*2048+ 567,   45*2048+ 568,   45*2048+ 569,   45*2048+ 570,    8*2048+ 571,   45*2048+ 572,   44*2048+ 573,   37*2048+ 574,    7*2048+ 575,   42*2048+ 576,   25*2048+ 577,   45*2048+ 578,   45*2048+ 579, 
  29*2048+ 580,   10*2048+ 581,   32*2048+ 582,   18*2048+ 583,   12*2048+ 584,   45*2048+ 585,   45*2048+ 586,   45*2048+ 587,   45*2048+ 588,   15*2048+ 589,   19*2048+ 590,   43*2048+ 591,    6*2048+ 592,   22*2048+ 593,   45*2048+ 594,   45*2048+ 595, 
  38*2048+ 596,   43*2048+ 597,   44*2048+ 598,   45*2048+ 599,   45*2048+ 600,   10*2048+ 601,   45*2048+ 602,   45*2048+ 603,   45*2048+ 604,   37*2048+ 605,   32*2048+ 606,    3*2048+ 607,   38*2048+ 608,   20*2048+ 609,   45*2048+ 610,   45*2048+ 611, 
  19*2048+ 685,   19*2048+ 686,   10*2048+ 687,    8*2048+ 688,   28*2048+ 689,    9*2048+ 690,   26*2048+ 691,   45*2048+ 692,   12*2048+ 693,   45*2048+ 694,   45*2048+ 695,   41*2048+ 696,   45*2048+ 697,   25*2048+ 698,   45*2048+ 699,   45*2048+ 700, 
   8*2048+ 701,   43*2048+ 702,   26*2048+ 703,   37*2048+ 704,   44*2048+ 705,   22*2048+ 706,   26*2048+ 707,   45*2048+ 708,   45*2048+ 709,   45*2048+ 710,    8*2048+ 711,   45*2048+ 712,   44*2048+ 713,   37*2048+ 714,   45*2048+ 715,   45*2048+ 716, 
  23*2048+ 717,   29*2048+ 718,   10*2048+ 719,   32*2048+ 720,   18*2048+ 721,   12*2048+ 722,   45*2048+ 723,   45*2048+ 724,   45*2048+ 725,   45*2048+ 726,   15*2048+ 727,   19*2048+ 728,   43*2048+ 729,    6*2048+ 730,   45*2048+ 731,   45*2048+ 732, 
  21*2048+ 733,   38*2048+ 734,   43*2048+ 735,   44*2048+ 736,   45*2048+ 737,   45*2048+ 738,   10*2048+ 739,   45*2048+ 740,   45*2048+ 741,   45*2048+ 742,   37*2048+ 743,   32*2048+ 744,    3*2048+ 745,   38*2048+ 746,   45*2048+ 747,   45*2048+ 748, 
  26*2048+ 822,   19*2048+ 823,   19*2048+ 824,   10*2048+ 825,    8*2048+ 826,   28*2048+ 827,    9*2048+ 828,   26*2048+ 829,   45*2048+ 830,   12*2048+ 831,   45*2048+ 832,   45*2048+ 833,   41*2048+ 834,   45*2048+ 835,   45*2048+ 836,   45*2048+ 837, 
  38*2048+ 838,    8*2048+ 839,   43*2048+ 840,   26*2048+ 841,   37*2048+ 842,   44*2048+ 843,   22*2048+ 844,   26*2048+ 845,   45*2048+ 846,   45*2048+ 847,   45*2048+ 848,    8*2048+ 849,   45*2048+ 850,   44*2048+ 851,   45*2048+ 852,   45*2048+ 853, 
  44*2048+ 854,    7*2048+ 855,   23*2048+ 856,   29*2048+ 857,   10*2048+ 858,   32*2048+ 859,   18*2048+ 860,   12*2048+ 861,   45*2048+ 862,   45*2048+ 863,   45*2048+ 864,   45*2048+ 865,   15*2048+ 866,   19*2048+ 867,   45*2048+ 868,   45*2048+ 869, 
  38*2048+ 870,   33*2048+ 871,    4*2048+ 872,   39*2048+ 873,   21*2048+ 874,   38*2048+ 875,   43*2048+ 876,   44*2048+ 877,   45*2048+ 878,   45*2048+ 879,   10*2048+ 880,   45*2048+ 881,   45*2048+ 882,   45*2048+ 883,   45*2048+ 884,   45*2048+ 885, 
  26*2048+ 959,   19*2048+ 960,   19*2048+ 961,   10*2048+ 962,    8*2048+ 963,   28*2048+ 964,    9*2048+ 965,   26*2048+ 966,   45*2048+ 967,   12*2048+ 968,   45*2048+ 969,   45*2048+ 970,   41*2048+ 971,   45*2048+ 972,   45*2048+ 973,   45*2048+ 974, 
  45*2048+ 975,   38*2048+ 976,    8*2048+ 977,   43*2048+ 978,   26*2048+ 979,   37*2048+ 980,   44*2048+ 981,   22*2048+ 982,   26*2048+ 983,   45*2048+ 984,   45*2048+ 985,   45*2048+ 986,    8*2048+ 987,   45*2048+ 988,   45*2048+ 989,   45*2048+ 990, 
  16*2048+ 991,   20*2048+ 992,   44*2048+ 993,    7*2048+ 994,   23*2048+ 995,   29*2048+ 996,   10*2048+ 997,   32*2048+ 998,   18*2048+ 999,   12*2048+1000,   45*2048+1001,   45*2048+1002,   45*2048+1003,   45*2048+1004,   45*2048+1005,   45*2048+1006, 
  38*2048+1007,   33*2048+1008,    4*2048+1009,   39*2048+1010,   21*2048+1011,   38*2048+1012,   43*2048+1013,   44*2048+1014,   45*2048+1015,   45*2048+1016,   10*2048+1017,   45*2048+1018,   45*2048+1019,   45*2048+1020,   45*2048+1021,   45*2048+1022, 
  45*2048+ 120,   45*2048+ 121,   33*2048+ 122,   45*2048+ 123,   45*2048+ 124,   45*2048+ 125,   37*2048+ 126,   30*2048+ 127,   36*2048+ 128,    6*2048+ 129,    7*2048+ 130,   42*2048+ 131,    0*2048+ 132,    5*2048+ 133,   25*2048+ 134,   45*2048+ 135,   45*2048+ 136, 
   7*2048+ 257,    8*2048+ 258,   43*2048+ 259,    1*2048+ 260,    6*2048+ 261,   26*2048+ 262,   45*2048+ 263,   45*2048+ 264,   33*2048+ 265,   45*2048+ 266,   45*2048+ 267,   45*2048+ 268,   37*2048+ 269,   30*2048+ 270,   36*2048+ 271,   45*2048+ 272,   45*2048+ 273, 
   7*2048+ 394,    8*2048+ 395,   43*2048+ 396,    1*2048+ 397,    6*2048+ 398,   26*2048+ 399,   45*2048+ 400,   45*2048+ 401,   33*2048+ 402,   45*2048+ 403,   45*2048+ 404,   45*2048+ 405,   37*2048+ 406,   30*2048+ 407,   36*2048+ 408,   45*2048+ 409,   45*2048+ 410, 
   7*2048+ 531,    8*2048+ 532,   43*2048+ 533,    1*2048+ 534,    6*2048+ 535,   26*2048+ 536,   45*2048+ 537,   45*2048+ 538,   33*2048+ 539,   45*2048+ 540,   45*2048+ 541,   45*2048+ 542,   37*2048+ 543,   30*2048+ 544,   36*2048+ 545,   45*2048+ 546,   45*2048+ 547, 
   7*2048+ 668,    8*2048+ 669,   43*2048+ 670,    1*2048+ 671,    6*2048+ 672,   26*2048+ 673,   45*2048+ 674,   45*2048+ 675,   33*2048+ 676,   45*2048+ 677,   45*2048+ 678,   45*2048+ 679,   37*2048+ 680,   30*2048+ 681,   36*2048+ 682,   45*2048+ 683,   45*2048+ 684, 
  37*2048+ 805,    7*2048+ 806,    8*2048+ 807,   43*2048+ 808,    1*2048+ 809,    6*2048+ 810,   26*2048+ 811,   45*2048+ 812,   45*2048+ 813,   33*2048+ 814,   45*2048+ 815,   45*2048+ 816,   45*2048+ 817,   37*2048+ 818,   30*2048+ 819,   45*2048+ 820,   45*2048+ 821, 
  38*2048+ 942,   31*2048+ 943,   37*2048+ 944,    7*2048+ 945,    8*2048+ 946,   43*2048+ 947,    1*2048+ 948,    6*2048+ 949,   26*2048+ 950,   45*2048+ 951,   45*2048+ 952,   33*2048+ 953,   45*2048+ 954,   45*2048+ 955,   45*2048+ 956,   45*2048+ 957,   45*2048+ 958, 
  38*2048+1079,   31*2048+1080,   37*2048+1081,    7*2048+1082,    8*2048+1083,   43*2048+1084,    1*2048+1085,    6*2048+1086,   26*2048+1087,   45*2048+1088,   45*2048+1089,   33*2048+1090,   45*2048+1091,   45*2048+1092,   45*2048+1093,   45*2048+1094,   45*2048+1095, 
  45*2048+  83,   45*2048+  84,   45*2048+  85,   45*2048+  86,   45*2048+  87,   35*2048+  88,   36*2048+  89,    1*2048+  90,    7*2048+  91,   20*2048+  92,   25*2048+  93,   18*2048+  94,   25*2048+  95,   27*2048+  96,   15*2048+  97,   39*2048+  98,   45*2048+  99,   45*2048+ 100, 
  40*2048+ 220,   45*2048+ 221,   45*2048+ 222,   45*2048+ 223,   45*2048+ 224,   45*2048+ 225,   35*2048+ 226,   36*2048+ 227,    1*2048+ 228,    7*2048+ 229,   20*2048+ 230,   25*2048+ 231,   18*2048+ 232,   25*2048+ 233,   27*2048+ 234,   15*2048+ 235,   45*2048+ 236,   45*2048+ 237, 
  40*2048+ 357,   45*2048+ 358,   45*2048+ 359,   45*2048+ 360,   45*2048+ 361,   45*2048+ 362,   35*2048+ 363,   36*2048+ 364,    1*2048+ 365,    7*2048+ 366,   20*2048+ 367,   25*2048+ 368,   18*2048+ 369,   25*2048+ 370,   27*2048+ 371,   15*2048+ 372,   45*2048+ 373,   45*2048+ 374, 
  26*2048+ 494,   28*2048+ 495,   16*2048+ 496,   40*2048+ 497,   45*2048+ 498,   45*2048+ 499,   45*2048+ 500,   45*2048+ 501,   45*2048+ 502,   35*2048+ 503,   36*2048+ 504,    1*2048+ 505,    7*2048+ 506,   20*2048+ 507,   25*2048+ 508,   18*2048+ 509,   45*2048+ 510,   45*2048+ 511, 
  19*2048+ 631,   26*2048+ 632,   28*2048+ 633,   16*2048+ 634,   40*2048+ 635,   45*2048+ 636,   45*2048+ 637,   45*2048+ 638,   45*2048+ 639,   45*2048+ 640,   35*2048+ 641,   36*2048+ 642,    1*2048+ 643,    7*2048+ 644,   20*2048+ 645,   25*2048+ 646,   45*2048+ 647,   45*2048+ 648, 
   8*2048+ 768,   21*2048+ 769,   26*2048+ 770,   19*2048+ 771,   26*2048+ 772,   28*2048+ 773,   16*2048+ 774,   40*2048+ 775,   45*2048+ 776,   45*2048+ 777,   45*2048+ 778,   45*2048+ 779,   45*2048+ 780,   35*2048+ 781,   36*2048+ 782,    1*2048+ 783,   45*2048+ 784,   45*2048+ 785, 
   2*2048+ 905,    8*2048+ 906,   21*2048+ 907,   26*2048+ 908,   19*2048+ 909,   26*2048+ 910,   28*2048+ 911,   16*2048+ 912,   40*2048+ 913,   45*2048+ 914,   45*2048+ 915,   45*2048+ 916,   45*2048+ 917,   45*2048+ 918,   35*2048+ 919,   36*2048+ 920,   45*2048+ 921,   45*2048+ 922, 
  37*2048+1042,    2*2048+1043,    8*2048+1044,   21*2048+1045,   26*2048+1046,   19*2048+1047,   26*2048+1048,   28*2048+1049,   16*2048+1050,   40*2048+1051,   45*2048+1052,   45*2048+1053,   45*2048+1054,   45*2048+1055,   45*2048+1056,   35*2048+1057,   45*2048+1058,   45*2048+1059, 
  45*2048+  64,   45*2048+  65,   30*2048+  66,   45*2048+  67,   45*2048+  68,   45*2048+  69,   44*2048+  70,   10*2048+  71,    8*2048+  72,   41*2048+  73,   41*2048+  74,   36*2048+  75,   29*2048+  76,    3*2048+  77,   30*2048+  78,   33*2048+  79,    5*2048+  80,   45*2048+  81,   45*2048+  82, 
  15*2048+ 101,   45*2048+ 102,   45*2048+ 103,   45*2048+ 104,   22*2048+ 105,   45*2048+ 106,   32*2048+ 107,   14*2048+ 108,   45*2048+ 109,   25*2048+ 110,   25*2048+ 111,    9*2048+ 112,   18*2048+ 113,   42*2048+ 114,   38*2048+ 115,    8*2048+ 116,   29*2048+ 117,   45*2048+ 118,   45*2048+ 119, 
  31*2048+ 201,   34*2048+ 202,    6*2048+ 203,   45*2048+ 204,   45*2048+ 205,   30*2048+ 206,   45*2048+ 207,   45*2048+ 208,   45*2048+ 209,   44*2048+ 210,   10*2048+ 211,    8*2048+ 212,   41*2048+ 213,   41*2048+ 214,   36*2048+ 215,   29*2048+ 216,    3*2048+ 217,   45*2048+ 218,   45*2048+ 219, 
  30*2048+ 238,   15*2048+ 239,   45*2048+ 240,   45*2048+ 241,   45*2048+ 242,   22*2048+ 243,   45*2048+ 244,   32*2048+ 245,   14*2048+ 246,   45*2048+ 247,   25*2048+ 248,   25*2048+ 249,    9*2048+ 250,   18*2048+ 251,   42*2048+ 252,   38*2048+ 253,    8*2048+ 254,   45*2048+ 255,   45*2048+ 256, 
  42*2048+ 338,   37*2048+ 339,   30*2048+ 340,    4*2048+ 341,   31*2048+ 342,   34*2048+ 343,    6*2048+ 344,   45*2048+ 345,   45*2048+ 346,   30*2048+ 347,   45*2048+ 348,   45*2048+ 349,   45*2048+ 350,   44*2048+ 351,   10*2048+ 352,    8*2048+ 353,   41*2048+ 354,   45*2048+ 355,   45*2048+ 356, 
   9*2048+ 375,   30*2048+ 376,   15*2048+ 377,   45*2048+ 378,   45*2048+ 379,   45*2048+ 380,   22*2048+ 381,   45*2048+ 382,   32*2048+ 383,   14*2048+ 384,   45*2048+ 385,   25*2048+ 386,   25*2048+ 387,    9*2048+ 388,   18*2048+ 389,   42*2048+ 390,   38*2048+ 391,   45*2048+ 392,   45*2048+ 393, 
  42*2048+ 475,   37*2048+ 476,   30*2048+ 477,    4*2048+ 478,   31*2048+ 479,   34*2048+ 480,    6*2048+ 481,   45*2048+ 482,   45*2048+ 483,   30*2048+ 484,   45*2048+ 485,   45*2048+ 486,   45*2048+ 487,   44*2048+ 488,   10*2048+ 489,    8*2048+ 490,   41*2048+ 491,   45*2048+ 492,   45*2048+ 493, 
  39*2048+ 512,    9*2048+ 513,   30*2048+ 514,   15*2048+ 515,   45*2048+ 516,   45*2048+ 517,   45*2048+ 518,   22*2048+ 519,   45*2048+ 520,   32*2048+ 521,   14*2048+ 522,   45*2048+ 523,   25*2048+ 524,   25*2048+ 525,    9*2048+ 526,   18*2048+ 527,   42*2048+ 528,   45*2048+ 529,   45*2048+ 530, 
  42*2048+ 612,   42*2048+ 613,   37*2048+ 614,   30*2048+ 615,    4*2048+ 616,   31*2048+ 617,   34*2048+ 618,    6*2048+ 619,   45*2048+ 620,   45*2048+ 621,   30*2048+ 622,   45*2048+ 623,   45*2048+ 624,   45*2048+ 625,   44*2048+ 626,   10*2048+ 627,    8*2048+ 628,   45*2048+ 629,   45*2048+ 630, 
  19*2048+ 649,   43*2048+ 650,   39*2048+ 651,    9*2048+ 652,   30*2048+ 653,   15*2048+ 654,   45*2048+ 655,   45*2048+ 656,   45*2048+ 657,   22*2048+ 658,   45*2048+ 659,   32*2048+ 660,   14*2048+ 661,   45*2048+ 662,   25*2048+ 663,   25*2048+ 664,    9*2048+ 665,   45*2048+ 666,   45*2048+ 667, 
   9*2048+ 749,   42*2048+ 750,   42*2048+ 751,   37*2048+ 752,   30*2048+ 753,    4*2048+ 754,   31*2048+ 755,   34*2048+ 756,    6*2048+ 757,   45*2048+ 758,   45*2048+ 759,   30*2048+ 760,   45*2048+ 761,   45*2048+ 762,   45*2048+ 763,   44*2048+ 764,   10*2048+ 765,   45*2048+ 766,   45*2048+ 767, 
  10*2048+ 786,   19*2048+ 787,   43*2048+ 788,   39*2048+ 789,    9*2048+ 790,   30*2048+ 791,   15*2048+ 792,   45*2048+ 793,   45*2048+ 794,   45*2048+ 795,   22*2048+ 796,   45*2048+ 797,   32*2048+ 798,   14*2048+ 799,   45*2048+ 800,   25*2048+ 801,   25*2048+ 802,   45*2048+ 803,   45*2048+ 804, 
  11*2048+ 886,    9*2048+ 887,   42*2048+ 888,   42*2048+ 889,   37*2048+ 890,   30*2048+ 891,    4*2048+ 892,   31*2048+ 893,   34*2048+ 894,    6*2048+ 895,   45*2048+ 896,   45*2048+ 897,   30*2048+ 898,   45*2048+ 899,   45*2048+ 900,   45*2048+ 901,   44*2048+ 902,   45*2048+ 903,   45*2048+ 904, 
  26*2048+ 923,   10*2048+ 924,   19*2048+ 925,   43*2048+ 926,   39*2048+ 927,    9*2048+ 928,   30*2048+ 929,   15*2048+ 930,   45*2048+ 931,   45*2048+ 932,   45*2048+ 933,   22*2048+ 934,   45*2048+ 935,   32*2048+ 936,   14*2048+ 937,   45*2048+ 938,   25*2048+ 939,   45*2048+ 940,   45*2048+ 941, 
  11*2048+1023,    9*2048+1024,   42*2048+1025,   42*2048+1026,   37*2048+1027,   30*2048+1028,    4*2048+1029,   31*2048+1030,   34*2048+1031,    6*2048+1032,   45*2048+1033,   45*2048+1034,   30*2048+1035,   45*2048+1036,   45*2048+1037,   45*2048+1038,   44*2048+1039,   45*2048+1040,   45*2048+1041, 
  26*2048+1060,   26*2048+1061,   10*2048+1062,   19*2048+1063,   43*2048+1064,   39*2048+1065,    9*2048+1066,   30*2048+1067,   15*2048+1068,   45*2048+1069,   45*2048+1070,   45*2048+1071,   22*2048+1072,   45*2048+1073,   32*2048+1074,   14*2048+1075,   45*2048+1076,   45*2048+1077,   45*2048+1078, 

  45*2048+   0,   45*2048+   1,   45*2048+   2,   45*2048+   3,   45*2048+   4,   21*2048+   5,   45*2048+   6,   45*2048+   7,   45*2048+   8,   20*2048+   9,   15*2048+  10,   24*2048+  11,   16*2048+  12,   16*2048+  13,    7*2048+  14,   15*2048+  15,   29*2048+  16,   35*2048+  17,    7*2048+  18,    7*2048+  19,   19*2048+  20,    8*2048+  21,   39*2048+  22,   24*2048+  23,   29*2048+  24,   45*2048+  25,   44*2048+  26, 
  45*2048+  27,   45*2048+  28,   45*2048+  29,   45*2048+  30,   45*2048+  31,   45*2048+  32,   45*2048+  33,   45*2048+  34,   31*2048+  35,   41*2048+  36,   41*2048+  37,   29*2048+  38,   32*2048+  39,    1*2048+  40,    2*2048+  41,   13*2048+  42,   34*2048+  43,    7*2048+  44,    8*2048+  45,   24*2048+  46,    5*2048+  47,   21*2048+  48,   10*2048+  49,   19*2048+  50,   13*2048+  51,   45*2048+  52,   45*2048+  53, 
  45*2048+  54,   33*2048+  55,   45*2048+  56,   45*2048+  57,   45*2048+  58,   45*2048+  59,   40*2048+  60,    2*2048+  61,   45*2048+  62,   45*2048+  63,   45*2048+  64,   27*2048+  65,    8*2048+  66,   35*2048+  67,   34*2048+  68,   32*2048+  69,   11*2048+  70,   25*2048+  71,   42*2048+  72,   28*2048+  73,   30*2048+  74,   27*2048+  75,   26*2048+  76,   15*2048+  77,   35*2048+  78,   45*2048+  79,   45*2048+  80, 
  45*2048+  81,   22*2048+  82,   45*2048+  83,   45*2048+  84,   10*2048+  85,   45*2048+  86,   12*2048+  87,   45*2048+  88,   45*2048+  89,   45*2048+  90,   45*2048+  91,    6*2048+  92,   37*2048+  93,   23*2048+  94,   24*2048+  95,    9*2048+  96,   32*2048+  97,    5*2048+  98,   17*2048+  99,   22*2048+ 100,    8*2048+ 101,   29*2048+ 102,   32*2048+ 103,   10*2048+ 104,   11*2048+ 105,   45*2048+ 106,   45*2048+ 107, 
  45*2048+ 108,   45*2048+ 109,    8*2048+ 110,   17*2048+ 111,   45*2048+ 112,   45*2048+ 113,   45*2048+ 114,    6*2048+ 115,   45*2048+ 116,   38*2048+ 117,   45*2048+ 118,   45*2048+ 119,   19*2048+ 120,   23*2048+ 121,   34*2048+ 122,   15*2048+ 123,   29*2048+ 124,   31*2048+ 125,    2*2048+ 126,   17*2048+ 127,   37*2048+ 128,   10*2048+ 129,   16*2048+ 130,   24*2048+ 131,   36*2048+ 132,   45*2048+ 133,   45*2048+ 134, 
  25*2048+ 135,   30*2048+ 136,   45*2048+ 137,   45*2048+ 138,   45*2048+ 139,   45*2048+ 140,   45*2048+ 141,   21*2048+ 142,   45*2048+ 143,   45*2048+ 144,   45*2048+ 145,   20*2048+ 146,   15*2048+ 147,   24*2048+ 148,   16*2048+ 149,   16*2048+ 150,    7*2048+ 151,   15*2048+ 152,   29*2048+ 153,   35*2048+ 154,    7*2048+ 155,    7*2048+ 156,   19*2048+ 157,    8*2048+ 158,   39*2048+ 159,   45*2048+ 160,   45*2048+ 161, 
  25*2048+ 162,    6*2048+ 163,   22*2048+ 164,   11*2048+ 165,   20*2048+ 166,   14*2048+ 167,   45*2048+ 168,   45*2048+ 169,   45*2048+ 170,   45*2048+ 171,   45*2048+ 172,   45*2048+ 173,   45*2048+ 174,   45*2048+ 175,   31*2048+ 176,   41*2048+ 177,   41*2048+ 178,   29*2048+ 179,   32*2048+ 180,    1*2048+ 181,    2*2048+ 182,   13*2048+ 183,   34*2048+ 184,    7*2048+ 185,    8*2048+ 186,   45*2048+ 187,   45*2048+ 188, 
  36*2048+ 189,   45*2048+ 190,   33*2048+ 191,   45*2048+ 192,   45*2048+ 193,   45*2048+ 194,   45*2048+ 195,   40*2048+ 196,    2*2048+ 197,   45*2048+ 198,   45*2048+ 199,   45*2048+ 200,   27*2048+ 201,    8*2048+ 202,   35*2048+ 203,   34*2048+ 204,   32*2048+ 205,   11*2048+ 206,   25*2048+ 207,   42*2048+ 208,   28*2048+ 209,   30*2048+ 210,   27*2048+ 211,   26*2048+ 212,   15*2048+ 213,   45*2048+ 214,   45*2048+ 215, 
  30*2048+ 216,   33*2048+ 217,   11*2048+ 218,   12*2048+ 219,   45*2048+ 220,   22*2048+ 221,   45*2048+ 222,   45*2048+ 223,   10*2048+ 224,   45*2048+ 225,   12*2048+ 226,   45*2048+ 227,   45*2048+ 228,   45*2048+ 229,   45*2048+ 230,    6*2048+ 231,   37*2048+ 232,   23*2048+ 233,   24*2048+ 234,    9*2048+ 235,   32*2048+ 236,    5*2048+ 237,   17*2048+ 238,   22*2048+ 239,    8*2048+ 240,   45*2048+ 241,   45*2048+ 242, 
  17*2048+ 243,   25*2048+ 244,   37*2048+ 245,   45*2048+ 246,   45*2048+ 247,    8*2048+ 248,   17*2048+ 249,   45*2048+ 250,   45*2048+ 251,   45*2048+ 252,    6*2048+ 253,   45*2048+ 254,   38*2048+ 255,   45*2048+ 256,   45*2048+ 257,   19*2048+ 258,   23*2048+ 259,   34*2048+ 260,   15*2048+ 261,   29*2048+ 262,   31*2048+ 263,    2*2048+ 264,   17*2048+ 265,   37*2048+ 266,   10*2048+ 267,   45*2048+ 268,   45*2048+ 269, 
   9*2048+ 270,   40*2048+ 271,   25*2048+ 272,   30*2048+ 273,   45*2048+ 274,   45*2048+ 275,   45*2048+ 276,   45*2048+ 277,   45*2048+ 278,   21*2048+ 279,   45*2048+ 280,   45*2048+ 281,   45*2048+ 282,   20*2048+ 283,   15*2048+ 284,   24*2048+ 285,   16*2048+ 286,   16*2048+ 287,    7*2048+ 288,   15*2048+ 289,   29*2048+ 290,   35*2048+ 291,    7*2048+ 292,    7*2048+ 293,   19*2048+ 294,   45*2048+ 295,   45*2048+ 296, 
   9*2048+ 297,   25*2048+ 298,    6*2048+ 299,   22*2048+ 300,   11*2048+ 301,   20*2048+ 302,   14*2048+ 303,   45*2048+ 304,   45*2048+ 305,   45*2048+ 306,   45*2048+ 307,   45*2048+ 308,   45*2048+ 309,   45*2048+ 310,   45*2048+ 311,   31*2048+ 312,   41*2048+ 313,   41*2048+ 314,   29*2048+ 315,   32*2048+ 316,    1*2048+ 317,    2*2048+ 318,   13*2048+ 319,   34*2048+ 320,    7*2048+ 321,   45*2048+ 322,   45*2048+ 323, 
  28*2048+ 324,   27*2048+ 325,   16*2048+ 326,   36*2048+ 327,   45*2048+ 328,   33*2048+ 329,   45*2048+ 330,   45*2048+ 331,   45*2048+ 332,   45*2048+ 333,   40*2048+ 334,    2*2048+ 335,   45*2048+ 336,   45*2048+ 337,   45*2048+ 338,   27*2048+ 339,    8*2048+ 340,   35*2048+ 341,   34*2048+ 342,   32*2048+ 343,   11*2048+ 344,   25*2048+ 345,   42*2048+ 346,   28*2048+ 347,   30*2048+ 348,   45*2048+ 349,   45*2048+ 350, 
   9*2048+ 351,   30*2048+ 352,   33*2048+ 353,   11*2048+ 354,   12*2048+ 355,   45*2048+ 356,   22*2048+ 357,   45*2048+ 358,   45*2048+ 359,   10*2048+ 360,   45*2048+ 361,   12*2048+ 362,   45*2048+ 363,   45*2048+ 364,   45*2048+ 365,   45*2048+ 366,    6*2048+ 367,   37*2048+ 368,   23*2048+ 369,   24*2048+ 370,    9*2048+ 371,   32*2048+ 372,    5*2048+ 373,   17*2048+ 374,   22*2048+ 375,   45*2048+ 376,   45*2048+ 377, 
  38*2048+ 378,   11*2048+ 379,   17*2048+ 380,   25*2048+ 381,   37*2048+ 382,   45*2048+ 383,   45*2048+ 384,    8*2048+ 385,   17*2048+ 386,   45*2048+ 387,   45*2048+ 388,   45*2048+ 389,    6*2048+ 390,   45*2048+ 391,   38*2048+ 392,   45*2048+ 393,   45*2048+ 394,   19*2048+ 395,   23*2048+ 396,   34*2048+ 397,   15*2048+ 398,   29*2048+ 399,   31*2048+ 400,    2*2048+ 401,   17*2048+ 402,   45*2048+ 403,   45*2048+ 404, 
   8*2048+ 405,   20*2048+ 406,    9*2048+ 407,   40*2048+ 408,   25*2048+ 409,   30*2048+ 410,   45*2048+ 411,   45*2048+ 412,   45*2048+ 413,   45*2048+ 414,   45*2048+ 415,   21*2048+ 416,   45*2048+ 417,   45*2048+ 418,   45*2048+ 419,   20*2048+ 420,   15*2048+ 421,   24*2048+ 422,   16*2048+ 423,   16*2048+ 424,    7*2048+ 425,   15*2048+ 426,   29*2048+ 427,   35*2048+ 428,    7*2048+ 429,   45*2048+ 430,   45*2048+ 431, 
   8*2048+ 432,    9*2048+ 433,   25*2048+ 434,    6*2048+ 435,   22*2048+ 436,   11*2048+ 437,   20*2048+ 438,   14*2048+ 439,   45*2048+ 440,   45*2048+ 441,   45*2048+ 442,   45*2048+ 443,   45*2048+ 444,   45*2048+ 445,   45*2048+ 446,   45*2048+ 447,   31*2048+ 448,   41*2048+ 449,   41*2048+ 450,   29*2048+ 451,   32*2048+ 452,    1*2048+ 453,    2*2048+ 454,   13*2048+ 455,   34*2048+ 456,   45*2048+ 457,   45*2048+ 458, 
  12*2048+ 459,   26*2048+ 460,   43*2048+ 461,   29*2048+ 462,   31*2048+ 463,   28*2048+ 464,   27*2048+ 465,   16*2048+ 466,   36*2048+ 467,   45*2048+ 468,   33*2048+ 469,   45*2048+ 470,   45*2048+ 471,   45*2048+ 472,   45*2048+ 473,   40*2048+ 474,    2*2048+ 475,   45*2048+ 476,   45*2048+ 477,   45*2048+ 478,   27*2048+ 479,    8*2048+ 480,   35*2048+ 481,   34*2048+ 482,   32*2048+ 483,   45*2048+ 484,   45*2048+ 485, 
   6*2048+ 486,   18*2048+ 487,   23*2048+ 488,    9*2048+ 489,   30*2048+ 490,   33*2048+ 491,   11*2048+ 492,   12*2048+ 493,   45*2048+ 494,   22*2048+ 495,   45*2048+ 496,   45*2048+ 497,   10*2048+ 498,   45*2048+ 499,   12*2048+ 500,   45*2048+ 501,   45*2048+ 502,   45*2048+ 503,   45*2048+ 504,    6*2048+ 505,   37*2048+ 506,   23*2048+ 507,   24*2048+ 508,    9*2048+ 509,   32*2048+ 510,   45*2048+ 511,   45*2048+ 512, 
  38*2048+ 513,   11*2048+ 514,   17*2048+ 515,   25*2048+ 516,   37*2048+ 517,   45*2048+ 518,   45*2048+ 519,    8*2048+ 520,   17*2048+ 521,   45*2048+ 522,   45*2048+ 523,   45*2048+ 524,    6*2048+ 525,   45*2048+ 526,   38*2048+ 527,   45*2048+ 528,   45*2048+ 529,   19*2048+ 530,   23*2048+ 531,   34*2048+ 532,   15*2048+ 533,   29*2048+ 534,   31*2048+ 535,    2*2048+ 536,   17*2048+ 537,   45*2048+ 538,   45*2048+ 539, 
   8*2048+ 540,    8*2048+ 541,   20*2048+ 542,    9*2048+ 543,   40*2048+ 544,   25*2048+ 545,   30*2048+ 546,   45*2048+ 547,   45*2048+ 548,   45*2048+ 549,   45*2048+ 550,   45*2048+ 551,   21*2048+ 552,   45*2048+ 553,   45*2048+ 554,   45*2048+ 555,   20*2048+ 556,   15*2048+ 557,   24*2048+ 558,   16*2048+ 559,   16*2048+ 560,    7*2048+ 561,   15*2048+ 562,   29*2048+ 563,   35*2048+ 564,   45*2048+ 565,   45*2048+ 566, 
   2*2048+ 567,    3*2048+ 568,   14*2048+ 569,   35*2048+ 570,    8*2048+ 571,    9*2048+ 572,   25*2048+ 573,    6*2048+ 574,   22*2048+ 575,   11*2048+ 576,   20*2048+ 577,   14*2048+ 578,   45*2048+ 579,   45*2048+ 580,   45*2048+ 581,   45*2048+ 582,   45*2048+ 583,   45*2048+ 584,   45*2048+ 585,   45*2048+ 586,   31*2048+ 587,   41*2048+ 588,   41*2048+ 589,   29*2048+ 590,   32*2048+ 591,   45*2048+ 592,   45*2048+ 593, 
  33*2048+ 594,   12*2048+ 595,   26*2048+ 596,   43*2048+ 597,   29*2048+ 598,   31*2048+ 599,   28*2048+ 600,   27*2048+ 601,   16*2048+ 602,   36*2048+ 603,   45*2048+ 604,   33*2048+ 605,   45*2048+ 606,   45*2048+ 607,   45*2048+ 608,   45*2048+ 609,   40*2048+ 610,    2*2048+ 611,   45*2048+ 612,   45*2048+ 613,   45*2048+ 614,   27*2048+ 615,    8*2048+ 616,   35*2048+ 617,   34*2048+ 618,   45*2048+ 619,   45*2048+ 620, 
   6*2048+ 621,   18*2048+ 622,   23*2048+ 623,    9*2048+ 624,   30*2048+ 625,   33*2048+ 626,   11*2048+ 627,   12*2048+ 628,   45*2048+ 629,   22*2048+ 630,   45*2048+ 631,   45*2048+ 632,   10*2048+ 633,   45*2048+ 634,   12*2048+ 635,   45*2048+ 636,   45*2048+ 637,   45*2048+ 638,   45*2048+ 639,    6*2048+ 640,   37*2048+ 641,   23*2048+ 642,   24*2048+ 643,    9*2048+ 644,   32*2048+ 645,   45*2048+ 646,   45*2048+ 647, 
  16*2048+ 648,   30*2048+ 649,   32*2048+ 650,    3*2048+ 651,   18*2048+ 652,   38*2048+ 653,   11*2048+ 654,   17*2048+ 655,   25*2048+ 656,   37*2048+ 657,   45*2048+ 658,   45*2048+ 659,    8*2048+ 660,   17*2048+ 661,   45*2048+ 662,   45*2048+ 663,   45*2048+ 664,    6*2048+ 665,   45*2048+ 666,   38*2048+ 667,   45*2048+ 668,   45*2048+ 669,   19*2048+ 670,   23*2048+ 671,   34*2048+ 672,   45*2048+ 673,   45*2048+ 674, 
  36*2048+ 675,    8*2048+ 676,    8*2048+ 677,   20*2048+ 678,    9*2048+ 679,   40*2048+ 680,   25*2048+ 681,   30*2048+ 682,   45*2048+ 683,   45*2048+ 684,   45*2048+ 685,   45*2048+ 686,   45*2048+ 687,   21*2048+ 688,   45*2048+ 689,   45*2048+ 690,   45*2048+ 691,   20*2048+ 692,   15*2048+ 693,   24*2048+ 694,   16*2048+ 695,   16*2048+ 696,    7*2048+ 697,   15*2048+ 698,   29*2048+ 699,   45*2048+ 700,   45*2048+ 701, 
  33*2048+ 702,    2*2048+ 703,    3*2048+ 704,   14*2048+ 705,   35*2048+ 706,    8*2048+ 707,    9*2048+ 708,   25*2048+ 709,    6*2048+ 710,   22*2048+ 711,   11*2048+ 712,   20*2048+ 713,   14*2048+ 714,   45*2048+ 715,   45*2048+ 716,   45*2048+ 717,   45*2048+ 718,   45*2048+ 719,   45*2048+ 720,   45*2048+ 721,   45*2048+ 722,   31*2048+ 723,   41*2048+ 724,   41*2048+ 725,   29*2048+ 726,   45*2048+ 727,   45*2048+ 728, 
  35*2048+ 729,   33*2048+ 730,   12*2048+ 731,   26*2048+ 732,   43*2048+ 733,   29*2048+ 734,   31*2048+ 735,   28*2048+ 736,   27*2048+ 737,   16*2048+ 738,   36*2048+ 739,   45*2048+ 740,   33*2048+ 741,   45*2048+ 742,   45*2048+ 743,   45*2048+ 744,   45*2048+ 745,   40*2048+ 746,    2*2048+ 747,   45*2048+ 748,   45*2048+ 749,   45*2048+ 750,   27*2048+ 751,    8*2048+ 752,   35*2048+ 753,   45*2048+ 754,   45*2048+ 755, 
  25*2048+ 756,   10*2048+ 757,   33*2048+ 758,    6*2048+ 759,   18*2048+ 760,   23*2048+ 761,    9*2048+ 762,   30*2048+ 763,   33*2048+ 764,   11*2048+ 765,   12*2048+ 766,   45*2048+ 767,   22*2048+ 768,   45*2048+ 769,   45*2048+ 770,   10*2048+ 771,   45*2048+ 772,   12*2048+ 773,   45*2048+ 774,   45*2048+ 775,   45*2048+ 776,   45*2048+ 777,    6*2048+ 778,   37*2048+ 779,   23*2048+ 780,   45*2048+ 781,   45*2048+ 782, 
  35*2048+ 783,   16*2048+ 784,   30*2048+ 785,   32*2048+ 786,    3*2048+ 787,   18*2048+ 788,   38*2048+ 789,   11*2048+ 790,   17*2048+ 791,   25*2048+ 792,   37*2048+ 793,   45*2048+ 794,   45*2048+ 795,    8*2048+ 796,   17*2048+ 797,   45*2048+ 798,   45*2048+ 799,   45*2048+ 800,    6*2048+ 801,   45*2048+ 802,   38*2048+ 803,   45*2048+ 804,   45*2048+ 805,   19*2048+ 806,   23*2048+ 807,   45*2048+ 808,   45*2048+ 809, 
  16*2048+ 810,   30*2048+ 811,   36*2048+ 812,    8*2048+ 813,    8*2048+ 814,   20*2048+ 815,    9*2048+ 816,   40*2048+ 817,   25*2048+ 818,   30*2048+ 819,   45*2048+ 820,   45*2048+ 821,   45*2048+ 822,   45*2048+ 823,   45*2048+ 824,   21*2048+ 825,   45*2048+ 826,   45*2048+ 827,   45*2048+ 828,   20*2048+ 829,   15*2048+ 830,   24*2048+ 831,   16*2048+ 832,   16*2048+ 833,    7*2048+ 834,   45*2048+ 835,   45*2048+ 836, 
  42*2048+ 837,   42*2048+ 838,   30*2048+ 839,   33*2048+ 840,    2*2048+ 841,    3*2048+ 842,   14*2048+ 843,   35*2048+ 844,    8*2048+ 845,    9*2048+ 846,   25*2048+ 847,    6*2048+ 848,   22*2048+ 849,   11*2048+ 850,   20*2048+ 851,   14*2048+ 852,   45*2048+ 853,   45*2048+ 854,   45*2048+ 855,   45*2048+ 856,   45*2048+ 857,   45*2048+ 858,   45*2048+ 859,   45*2048+ 860,   31*2048+ 861,   45*2048+ 862,   45*2048+ 863, 
  28*2048+ 864,    9*2048+ 865,   36*2048+ 866,   35*2048+ 867,   33*2048+ 868,   12*2048+ 869,   26*2048+ 870,   43*2048+ 871,   29*2048+ 872,   31*2048+ 873,   28*2048+ 874,   27*2048+ 875,   16*2048+ 876,   36*2048+ 877,   45*2048+ 878,   33*2048+ 879,   45*2048+ 880,   45*2048+ 881,   45*2048+ 882,   45*2048+ 883,   40*2048+ 884,    2*2048+ 885,   45*2048+ 886,   45*2048+ 887,   45*2048+ 888,   45*2048+ 889,   45*2048+ 890, 
  24*2048+ 891,   25*2048+ 892,   10*2048+ 893,   33*2048+ 894,    6*2048+ 895,   18*2048+ 896,   23*2048+ 897,    9*2048+ 898,   30*2048+ 899,   33*2048+ 900,   11*2048+ 901,   12*2048+ 902,   45*2048+ 903,   22*2048+ 904,   45*2048+ 905,   45*2048+ 906,   10*2048+ 907,   45*2048+ 908,   12*2048+ 909,   45*2048+ 910,   45*2048+ 911,   45*2048+ 912,   45*2048+ 913,    6*2048+ 914,   37*2048+ 915,   45*2048+ 916,   45*2048+ 917, 
  24*2048+ 918,   35*2048+ 919,   16*2048+ 920,   30*2048+ 921,   32*2048+ 922,    3*2048+ 923,   18*2048+ 924,   38*2048+ 925,   11*2048+ 926,   17*2048+ 927,   25*2048+ 928,   37*2048+ 929,   45*2048+ 930,   45*2048+ 931,    8*2048+ 932,   17*2048+ 933,   45*2048+ 934,   45*2048+ 935,   45*2048+ 936,    6*2048+ 937,   45*2048+ 938,   38*2048+ 939,   45*2048+ 940,   45*2048+ 941,   19*2048+ 942,   45*2048+ 943,   45*2048+ 944, 
  16*2048+ 945,   25*2048+ 946,   17*2048+ 947,   17*2048+ 948,    8*2048+ 949,   16*2048+ 950,   30*2048+ 951,   36*2048+ 952,    8*2048+ 953,    8*2048+ 954,   20*2048+ 955,    9*2048+ 956,   40*2048+ 957,   25*2048+ 958,   30*2048+ 959,   45*2048+ 960,   45*2048+ 961,   45*2048+ 962,   45*2048+ 963,   45*2048+ 964,   21*2048+ 965,   45*2048+ 966,   45*2048+ 967,   45*2048+ 968,   20*2048+ 969,   45*2048+ 970,   45*2048+ 971, 
  32*2048+ 972,   42*2048+ 973,   42*2048+ 974,   30*2048+ 975,   33*2048+ 976,    2*2048+ 977,    3*2048+ 978,   14*2048+ 979,   35*2048+ 980,    8*2048+ 981,    9*2048+ 982,   25*2048+ 983,    6*2048+ 984,   22*2048+ 985,   11*2048+ 986,   20*2048+ 987,   14*2048+ 988,   45*2048+ 989,   45*2048+ 990,   45*2048+ 991,   45*2048+ 992,   45*2048+ 993,   45*2048+ 994,   45*2048+ 995,   45*2048+ 996,   45*2048+ 997,   45*2048+ 998, 
  28*2048+ 999,    9*2048+1000,   36*2048+1001,   35*2048+1002,   33*2048+1003,   12*2048+1004,   26*2048+1005,   43*2048+1006,   29*2048+1007,   31*2048+1008,   28*2048+1009,   27*2048+1010,   16*2048+1011,   36*2048+1012,   45*2048+1013,   33*2048+1014,   45*2048+1015,   45*2048+1016,   45*2048+1017,   45*2048+1018,   40*2048+1019,    2*2048+1020,   45*2048+1021,   45*2048+1022,   45*2048+1023,   45*2048+1024,   45*2048+1025, 
   7*2048+1026,   38*2048+1027,   24*2048+1028,   25*2048+1029,   10*2048+1030,   33*2048+1031,    6*2048+1032,   18*2048+1033,   23*2048+1034,    9*2048+1035,   30*2048+1036,   33*2048+1037,   11*2048+1038,   12*2048+1039,   45*2048+1040,   22*2048+1041,   45*2048+1042,   45*2048+1043,   10*2048+1044,   45*2048+1045,   12*2048+1046,   45*2048+1047,   45*2048+1048,   45*2048+1049,   45*2048+1050,   45*2048+1051,   45*2048+1052, 
  20*2048+1053,   24*2048+1054,   35*2048+1055,   16*2048+1056,   30*2048+1057,   32*2048+1058,    3*2048+1059,   18*2048+1060,   38*2048+1061,   11*2048+1062,   17*2048+1063,   25*2048+1064,   37*2048+1065,   45*2048+1066,   45*2048+1067,    8*2048+1068,   17*2048+1069,   45*2048+1070,   45*2048+1071,   45*2048+1072,    6*2048+1073,   45*2048+1074,   38*2048+1075,   45*2048+1076,   45*2048+1077,   45*2048+1078,   45*2048+1079);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if RdAddr < ROM'length then
				Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , Do'length );
			end if;
		end if;
	end process;

end Behavioral;