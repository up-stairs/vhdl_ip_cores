LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VNP_Output_Edge_Memory is
	Port (
		clk			: in  std_logic;

		RdAddr		: in  std_logic_vector(13 downto 0);
		Do			: out std_logic_vector(16 downto 0)
	);
end VNP_Output_Edge_Memory;

architecture Behavioral of VNP_Output_Edge_Memory is
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 15272-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
   0*2048+   2,    0*2048+   6,    0*2048+1152,
   0*2048+   7,    0*2048+  10,    0*2048+1153,
   0*2048+  11,    0*2048+  14,    0*2048+1154,
   0*2048+  15,    0*2048+  18,    0*2048+1155,
   0*2048+  19,    0*2048+  22,    0*2048+1156,
   0*2048+  23,    0*2048+  25,    0*2048+1157,
   0*2048+  26,    0*2048+  29,    0*2048+1158,
   0*2048+  30,    0*2048+  33,    0*2048+1159,
   0*2048+  34,    0*2048+  37,    0*2048+1160,
   0*2048+  38,    0*2048+  41,    0*2048+1161,
   0*2048+  42,    0*2048+  45,    0*2048+1162,
   0*2048+  46,    0*2048+  49,    0*2048+1163,
   0*2048+  50,    0*2048+  52,    0*2048+1164,
   0*2048+  53,    0*2048+  55,    0*2048+1165,
   0*2048+  56,    0*2048+  58,    0*2048+1166,
   0*2048+  59,    0*2048+  62,    0*2048+1167,
   0*2048+  63,    0*2048+  66,    0*2048+1168,
   0*2048+  67,    0*2048+  70,    0*2048+1169,
   0*2048+  71,    0*2048+  74,    0*2048+1170,
   0*2048+  75,    0*2048+  77,    0*2048+1171,
   0*2048+  78,    0*2048+  81,    0*2048+1172,
   0*2048+  82,    0*2048+  85,    0*2048+1173,
   0*2048+  86,    0*2048+  89,    0*2048+1174,
   0*2048+  90,    0*2048+  93,    0*2048+1175,
   0*2048+  94,    0*2048+  97,    0*2048+1176,
   0*2048+  98,    0*2048+ 100,    0*2048+1177,
   0*2048+ 101,    0*2048+ 103,    0*2048+1178,
   0*2048+ 104,    0*2048+ 106,    0*2048+1179,
   0*2048+ 107,    0*2048+ 110,    0*2048+1180,
   0*2048+ 111,    0*2048+ 113,    0*2048+1181,
   0*2048+ 114,    0*2048+ 117,    0*2048+1182,
   0*2048+ 118,    0*2048+ 121,    0*2048+1183,
   0*2048+ 122,    0*2048+ 125,    0*2048+1184,
   0*2048+ 126,    0*2048+ 129,    0*2048+1185,
   0*2048+ 130,    0*2048+ 133,    0*2048+1186,
   0*2048+ 134,    0*2048+ 137,    0*2048+1187,
   0*2048+ 138,    0*2048+ 141,    0*2048+1188,
   0*2048+ 142,    0*2048+ 145,    0*2048+1189,
   0*2048+ 146,    0*2048+ 149,    0*2048+1190,
   0*2048+ 150,    0*2048+ 153,    0*2048+1191,
   0*2048+ 154,    0*2048+ 157,    0*2048+1192,
   0*2048+ 158,    0*2048+ 160,    0*2048+1193,
   0*2048+ 161,    0*2048+ 164,    0*2048+1194,
   0*2048+ 165,    0*2048+ 168,    0*2048+1195,
   0*2048+ 169,    0*2048+ 172,    0*2048+1196,
   0*2048+ 173,    0*2048+ 176,    0*2048+1197,
   0*2048+ 177,    0*2048+ 180,    0*2048+1198,
   0*2048+ 181,    0*2048+ 184,    0*2048+1199,
   0*2048+ 185,    0*2048+ 187,    0*2048+1200,
   0*2048+ 188,    0*2048+ 190,    0*2048+1201,
   0*2048+ 191,    0*2048+ 193,    0*2048+1202,
   0*2048+ 194,    0*2048+ 197,    0*2048+1203,
   0*2048+ 198,    0*2048+ 201,    0*2048+1204,
   0*2048+ 202,    0*2048+ 205,    0*2048+1205,
   0*2048+ 206,    0*2048+ 209,    0*2048+1206,
   0*2048+ 210,    0*2048+ 212,    0*2048+1207,
   0*2048+ 213,    0*2048+ 216,    0*2048+1208,
   0*2048+ 217,    0*2048+ 220,    0*2048+1209,
   0*2048+ 221,    0*2048+ 224,    0*2048+1210,
   0*2048+ 225,    0*2048+ 228,    0*2048+1211,
   0*2048+ 229,    0*2048+ 232,    0*2048+1212,
   0*2048+ 233,    0*2048+ 235,    0*2048+1213,
   0*2048+ 236,    0*2048+ 238,    0*2048+1214,
   0*2048+ 239,    0*2048+ 241,    0*2048+1215,
   0*2048+ 242,    0*2048+ 245,    0*2048+1216,
   0*2048+ 246,    0*2048+ 248,    0*2048+1217,
   0*2048+ 249,    0*2048+ 252,    0*2048+1218,
   0*2048+ 253,    0*2048+ 256,    0*2048+1219,
   0*2048+ 257,    0*2048+ 260,    0*2048+1220,
   0*2048+ 261,    0*2048+ 264,    0*2048+1221,
   0*2048+ 265,    0*2048+ 268,    0*2048+1222,
   0*2048+ 269,    0*2048+ 272,    0*2048+1223,
   0*2048+ 273,    0*2048+ 276,    0*2048+1224,
   0*2048+ 277,    0*2048+ 280,    0*2048+1225,
   0*2048+ 281,    0*2048+ 284,    0*2048+1226,
   0*2048+ 285,    0*2048+ 288,    0*2048+1227,
   0*2048+ 289,    0*2048+ 292,    0*2048+1228,
   0*2048+ 293,    0*2048+ 295,    0*2048+1229,
   0*2048+ 296,    0*2048+ 299,    0*2048+1230,
   0*2048+ 300,    0*2048+ 303,    0*2048+1231,
   0*2048+ 304,    0*2048+ 307,    0*2048+1232,
   0*2048+ 308,    0*2048+ 311,    0*2048+1233,
   0*2048+ 312,    0*2048+ 315,    0*2048+1234,
   0*2048+ 316,    0*2048+ 319,    0*2048+1235,
   0*2048+ 320,    0*2048+ 322,    0*2048+1236,
   0*2048+ 323,    0*2048+ 325,    0*2048+1237,
   0*2048+ 326,    0*2048+ 328,    0*2048+1238,
   0*2048+ 329,    0*2048+ 332,    0*2048+1239,
   0*2048+ 333,    0*2048+ 336,    0*2048+1240,
   0*2048+ 337,    0*2048+ 340,    0*2048+1241,
   0*2048+ 341,    0*2048+ 344,    0*2048+1242,
   0*2048+ 345,    0*2048+ 347,    0*2048+1243,
   0*2048+ 348,    0*2048+ 351,    0*2048+1244,
   0*2048+ 352,    0*2048+ 355,    0*2048+1245,
   0*2048+ 356,    0*2048+ 359,    0*2048+1246,
   0*2048+ 360,    0*2048+ 363,    0*2048+1247,
   0*2048+ 364,    0*2048+ 367,    0*2048+1248,
   0*2048+ 368,    0*2048+ 370,    0*2048+1249,
   0*2048+ 371,    0*2048+ 373,    0*2048+1250,
   0*2048+ 374,    0*2048+ 376,    0*2048+1251,
   0*2048+ 377,    0*2048+ 380,    0*2048+1252,
   0*2048+ 381,    0*2048+ 383,    0*2048+1253,
   0*2048+ 384,    0*2048+ 387,    0*2048+1254,
   0*2048+ 388,    0*2048+ 391,    0*2048+1255,
   0*2048+ 392,    0*2048+ 395,    0*2048+1256,
   0*2048+ 396,    0*2048+ 399,    0*2048+1257,
   0*2048+ 400,    0*2048+ 403,    0*2048+1258,
   0*2048+ 404,    0*2048+ 407,    0*2048+1259,
   0*2048+ 408,    0*2048+ 411,    0*2048+1260,
   0*2048+ 412,    0*2048+ 415,    0*2048+1261,
   0*2048+ 416,    0*2048+ 419,    0*2048+1262,
   0*2048+ 420,    0*2048+ 423,    0*2048+1263,
   0*2048+ 424,    0*2048+ 427,    0*2048+1264,
   0*2048+ 428,    0*2048+ 430,    0*2048+1265,
   0*2048+ 431,    0*2048+ 434,    0*2048+1266,
   0*2048+ 435,    0*2048+ 438,    0*2048+1267,
   0*2048+ 439,    0*2048+ 442,    0*2048+1268,
   0*2048+ 443,    0*2048+ 446,    0*2048+1269,
   0*2048+ 447,    0*2048+ 450,    0*2048+1270,
   0*2048+ 451,    0*2048+ 454,    0*2048+1271,
   0*2048+ 455,    0*2048+ 457,    0*2048+1272,
   0*2048+ 458,    0*2048+ 460,    0*2048+1273,
   0*2048+ 461,    0*2048+ 463,    0*2048+1274,
   0*2048+ 464,    0*2048+ 467,    0*2048+1275,
   0*2048+ 468,    0*2048+ 471,    0*2048+1276,
   0*2048+ 472,    0*2048+ 475,    0*2048+1277,
   0*2048+ 476,    0*2048+ 479,    0*2048+1278,
   0*2048+ 480,    0*2048+ 482,    0*2048+1279,
   0*2048+ 483,    0*2048+ 486,    0*2048+1280,
   0*2048+ 487,    0*2048+ 490,    0*2048+1281,
   0*2048+ 491,    0*2048+ 494,    0*2048+1282,
   0*2048+ 495,    0*2048+ 498,    0*2048+1283,
   0*2048+ 499,    0*2048+ 502,    0*2048+1284,
   0*2048+ 503,    0*2048+ 505,    0*2048+1285,
   0*2048+ 506,    0*2048+ 508,    0*2048+1286,
   0*2048+ 509,    0*2048+ 511,    0*2048+1287,
   0*2048+ 512,    0*2048+ 515,    0*2048+1288,
   0*2048+ 516,    0*2048+ 518,    0*2048+1289,
   0*2048+ 519,    0*2048+ 522,    0*2048+1290,
   0*2048+ 523,    0*2048+ 526,    0*2048+1291,
   0*2048+ 527,    0*2048+ 530,    0*2048+1292,
   0*2048+ 531,    0*2048+ 534,    0*2048+1293,
   0*2048+ 535,    0*2048+ 538,    0*2048+1294,
   0*2048+ 539,    0*2048+ 542,    0*2048+1295,
   0*2048+ 543,    0*2048+ 546,    0*2048+1296,
   0*2048+ 547,    0*2048+ 550,    0*2048+1297,
   0*2048+ 551,    0*2048+ 554,    0*2048+1298,
   0*2048+ 555,    0*2048+ 558,    0*2048+1299,
   0*2048+ 559,    0*2048+ 562,    0*2048+1300,
   0*2048+ 563,    0*2048+ 565,    0*2048+1301,
   0*2048+ 566,    0*2048+ 569,    0*2048+1302,
   0*2048+ 570,    0*2048+ 573,    0*2048+1303,
   0*2048+ 574,    0*2048+ 577,    0*2048+1304,
   0*2048+ 578,    0*2048+ 581,    0*2048+1305,
   0*2048+ 582,    0*2048+ 585,    0*2048+1306,
   0*2048+ 586,    0*2048+ 589,    0*2048+1307,
   0*2048+ 590,    0*2048+ 592,    0*2048+1308,
   0*2048+ 593,    0*2048+ 595,    0*2048+1309,
   0*2048+ 596,    0*2048+ 598,    0*2048+1310,
   0*2048+ 599,    0*2048+ 602,    0*2048+1311,
   0*2048+ 603,    0*2048+ 606,    0*2048+1312,
   0*2048+ 607,    0*2048+ 610,    0*2048+1313,
   0*2048+ 611,    0*2048+ 614,    0*2048+1314,
   0*2048+ 615,    0*2048+ 617,    0*2048+1315,
   0*2048+ 618,    0*2048+ 621,    0*2048+1316,
   0*2048+ 622,    0*2048+ 625,    0*2048+1317,
   0*2048+ 626,    0*2048+ 629,    0*2048+1318,
   0*2048+ 630,    0*2048+ 633,    0*2048+1319,
   0*2048+ 634,    0*2048+ 637,    0*2048+1320,
   0*2048+ 638,    0*2048+ 640,    0*2048+1321,
   0*2048+ 641,    0*2048+ 643,    0*2048+1322,
   0*2048+ 644,    0*2048+ 646,    0*2048+1323,
   0*2048+ 647,    0*2048+ 650,    0*2048+1324,
   0*2048+ 651,    0*2048+ 653,    0*2048+1325,
   0*2048+ 654,    0*2048+ 657,    0*2048+1326,
   0*2048+ 658,    0*2048+ 661,    0*2048+1327,
   0*2048+ 662,    0*2048+ 665,    0*2048+1328,
   0*2048+ 666,    0*2048+ 669,    0*2048+1329,
   0*2048+ 670,    0*2048+ 673,    0*2048+1330,
   0*2048+ 674,    0*2048+ 677,    0*2048+1331,
   0*2048+ 678,    0*2048+ 681,    0*2048+1332,
   0*2048+ 682,    0*2048+ 685,    0*2048+1333,
   0*2048+ 686,    0*2048+ 689,    0*2048+1334,
   0*2048+ 690,    0*2048+ 693,    0*2048+1335,
   0*2048+ 694,    0*2048+ 697,    0*2048+1336,
   0*2048+ 698,    0*2048+ 700,    0*2048+1337,
   0*2048+ 701,    0*2048+ 704,    0*2048+1338,
   0*2048+ 705,    0*2048+ 708,    0*2048+1339,
   0*2048+ 709,    0*2048+ 712,    0*2048+1340,
   0*2048+ 713,    0*2048+ 716,    0*2048+1341,
   0*2048+ 717,    0*2048+ 720,    0*2048+1342,
   0*2048+ 721,    0*2048+ 724,    0*2048+1343,
   0*2048+ 725,    0*2048+ 727,    0*2048+1344,
   0*2048+ 728,    0*2048+ 730,    0*2048+1345,
   0*2048+ 731,    0*2048+ 733,    0*2048+1346,
   0*2048+ 734,    0*2048+ 737,    0*2048+1347,
   0*2048+ 738,    0*2048+ 741,    0*2048+1348,
   0*2048+ 742,    0*2048+ 745,    0*2048+1349,
   0*2048+ 746,    0*2048+ 749,    0*2048+1350,
   0*2048+ 750,    0*2048+ 752,    0*2048+1351,
   0*2048+ 753,    0*2048+ 756,    0*2048+1352,
   0*2048+ 757,    0*2048+ 760,    0*2048+1353,
   0*2048+ 761,    0*2048+ 764,    0*2048+1354,
   0*2048+ 765,    0*2048+ 768,    0*2048+1355,
   0*2048+ 769,    0*2048+ 772,    0*2048+1356,
   0*2048+ 773,    0*2048+ 775,    0*2048+1357,
   0*2048+ 776,    0*2048+ 778,    0*2048+1358,
   0*2048+ 779,    0*2048+ 781,    0*2048+1359,
   0*2048+ 782,    0*2048+ 785,    0*2048+1360,
   0*2048+ 786,    0*2048+ 788,    0*2048+1361,
   0*2048+ 789,    0*2048+ 792,    0*2048+1362,
   0*2048+ 793,    0*2048+ 796,    0*2048+1363,
   0*2048+ 797,    0*2048+ 800,    0*2048+1364,
   0*2048+ 801,    0*2048+ 804,    0*2048+1365,
   0*2048+ 805,    0*2048+ 808,    0*2048+1366,
   0*2048+ 809,    0*2048+ 812,    0*2048+1367,
   0*2048+ 813,    0*2048+ 816,    0*2048+1368,
   0*2048+ 817,    0*2048+ 820,    0*2048+1369,
   0*2048+ 821,    0*2048+ 824,    0*2048+1370,
   0*2048+ 825,    0*2048+ 828,    0*2048+1371,
   0*2048+ 829,    0*2048+ 832,    0*2048+1372,
   0*2048+ 833,    0*2048+ 835,    0*2048+1373,
   0*2048+ 836,    0*2048+ 839,    0*2048+1374,
   0*2048+ 840,    0*2048+ 843,    0*2048+1375,
   0*2048+ 844,    0*2048+ 847,    0*2048+1376,
   0*2048+ 848,    0*2048+ 851,    0*2048+1377,
   0*2048+ 852,    0*2048+ 855,    0*2048+1378,
   0*2048+ 856,    0*2048+ 859,    0*2048+1379,
   0*2048+ 860,    0*2048+ 862,    0*2048+1380,
   0*2048+ 863,    0*2048+ 865,    0*2048+1381,
   0*2048+ 866,    0*2048+ 868,    0*2048+1382,
   0*2048+ 869,    0*2048+ 872,    0*2048+1383,
   0*2048+ 873,    0*2048+ 876,    0*2048+1384,
   0*2048+ 877,    0*2048+ 880,    0*2048+1385,
   0*2048+ 881,    0*2048+ 884,    0*2048+1386,
   0*2048+ 885,    0*2048+ 887,    0*2048+1387,
   0*2048+ 888,    0*2048+ 891,    0*2048+1388,
   0*2048+ 892,    0*2048+ 895,    0*2048+1389,
   0*2048+ 896,    0*2048+ 899,    0*2048+1390,
   0*2048+ 900,    0*2048+ 903,    0*2048+1391,
   0*2048+ 904,    0*2048+ 907,    0*2048+1392,
   0*2048+ 908,    0*2048+ 910,    0*2048+1393,
   0*2048+ 911,    0*2048+ 913,    0*2048+1394,
   0*2048+ 914,    0*2048+ 916,    0*2048+1395,
   0*2048+ 917,    0*2048+ 920,    0*2048+1396,
   0*2048+ 921,    0*2048+ 923,    0*2048+1397,
   0*2048+ 924,    0*2048+ 927,    0*2048+1398,
   0*2048+ 928,    0*2048+ 931,    0*2048+1399,
   0*2048+ 932,    0*2048+ 935,    0*2048+1400,
   0*2048+ 936,    0*2048+ 939,    0*2048+1401,
   0*2048+ 940,    0*2048+ 943,    0*2048+1402,
   0*2048+ 944,    0*2048+ 947,    0*2048+1403,
   0*2048+ 948,    0*2048+ 951,    0*2048+1404,
   0*2048+ 952,    0*2048+ 955,    0*2048+1405,
   0*2048+ 956,    0*2048+ 959,    0*2048+1406,
   0*2048+ 960,    0*2048+ 963,    0*2048+1407,
   0*2048+ 964,    0*2048+ 967,    0*2048+1408,
   0*2048+ 968,    0*2048+ 970,    0*2048+1409,
   0*2048+ 971,    0*2048+ 974,    0*2048+1410,
   0*2048+ 975,    0*2048+ 978,    0*2048+1411,
   0*2048+ 979,    0*2048+ 982,    0*2048+1412,
   0*2048+ 983,    0*2048+ 986,    0*2048+1413,
   0*2048+ 987,    0*2048+ 990,    0*2048+1414,
   0*2048+ 991,    0*2048+ 994,    0*2048+1415,
   0*2048+ 995,    0*2048+ 997,    0*2048+1416,
   0*2048+ 998,    0*2048+1000,    0*2048+1417,
   0*2048+1001,    0*2048+1003,    0*2048+1418,
   0*2048+1004,    0*2048+1007,    0*2048+1419,
   0*2048+1008,    0*2048+1011,    0*2048+1420,
   0*2048+1012,    0*2048+1015,    0*2048+1421,
   0*2048+1016,    0*2048+1019,    0*2048+1422,
   0*2048+1020,    0*2048+1022,    0*2048+1423,
   0*2048+1023,    0*2048+1026,    0*2048+1424,
   0*2048+1027,    0*2048+1030,    0*2048+1425,
   0*2048+1031,    0*2048+1034,    0*2048+1426,
   0*2048+1035,    0*2048+1038,    0*2048+1427,
   0*2048+1039,    0*2048+1042,    0*2048+1428,
   0*2048+1043,    0*2048+1045,    0*2048+1429,
   0*2048+1046,    0*2048+1048,    0*2048+1430,
   0*2048+1049,    0*2048+1051,    0*2048+1431,
   0*2048+1052,    0*2048+1055,    0*2048+1432,
   0*2048+1056,    0*2048+1058,    0*2048+1433,
   0*2048+1059,    0*2048+1062,    0*2048+1434,
   0*2048+1063,    0*2048+1066,    0*2048+1435,
   0*2048+1067,    0*2048+1070,    0*2048+1436,
   0*2048+1071,    0*2048+1074,    0*2048+1437,
   0*2048+1075,    0*2048+1078,    0*2048+1438,
   1*2048+   3,    0*2048+1079,    0*2048+1439,
  27*2048+ 254,   37*2048+ 440,   10*2048+ 748,    0*2048+1084,
  37*2048+ 743,   11*2048+ 814,   19*2048+1032,    0*2048+1085,
  42*2048+ 398,   41*2048+ 758,    4*2048+ 780,    0*2048+1086,
   8*2048+ 148,   21*2048+ 528,   14*2048+ 783,    0*2048+1087,
  34*2048+ 182,   44*2048+ 203,   17*2048+ 305,    0*2048+1088,
  27*2048+ 389,   37*2048+ 575,   10*2048+ 883,    0*2048+1093,
  20*2048+  87,   37*2048+ 878,   11*2048+ 949,    0*2048+1094,
  42*2048+ 533,   41*2048+ 893,    4*2048+ 915,    0*2048+1095,
   8*2048+ 283,   21*2048+ 663,   14*2048+ 918,    0*2048+1096,
  34*2048+ 317,   44*2048+ 338,   17*2048+ 441,    0*2048+1097,
  27*2048+ 524,   37*2048+ 710,   10*2048+1018,    0*2048+1102,
  12*2048+   4,   20*2048+ 222,   37*2048+1013,    0*2048+1103,
  42*2048+ 668,   41*2048+1028,    4*2048+1050,    0*2048+1104,
   8*2048+ 418,   21*2048+ 798,   14*2048+1053,    0*2048+1105,
  34*2048+ 452,   44*2048+ 473,   17*2048+ 576,    0*2048+1106,
  11*2048+  73,   27*2048+ 660,   37*2048+ 845,    0*2048+1111,
  38*2048+  68,   12*2048+ 139,   20*2048+ 358,    0*2048+1112,
  42*2048+  83,    5*2048+ 105,   42*2048+ 803,    0*2048+1113,
  15*2048+ 108,    8*2048+ 553,   21*2048+ 933,    0*2048+1114,
  34*2048+ 587,   44*2048+ 608,   17*2048+ 711,    0*2048+1115,
  11*2048+ 208,   27*2048+ 795,   37*2048+ 980,    0*2048+1120,
  38*2048+ 204,   12*2048+ 274,   20*2048+ 493,    0*2048+1121,
  42*2048+ 218,    5*2048+ 240,   42*2048+ 938,    0*2048+1122,
  15*2048+ 243,    8*2048+ 688,   21*2048+1068,    0*2048+1123,
  34*2048+ 722,   44*2048+ 744,   17*2048+ 846,    0*2048+1124,
  38*2048+  35,   11*2048+ 343,   27*2048+ 930,    0*2048+1129,
  38*2048+ 339,   12*2048+ 409,   20*2048+ 628,    0*2048+1130,
  42*2048+ 353,    5*2048+ 375,   42*2048+1073,    0*2048+1131,
  22*2048+ 123,   15*2048+ 378,    8*2048+ 823,    0*2048+1132,
  34*2048+ 857,   44*2048+ 879,   17*2048+ 981,    0*2048+1133,
  38*2048+ 170,   11*2048+ 478,   27*2048+1065,    0*2048+1138,
  38*2048+ 474,   12*2048+ 544,   20*2048+ 763,    0*2048+1139,
  43*2048+ 128,   42*2048+ 488,    5*2048+ 510,    0*2048+1140,
  22*2048+ 259,   15*2048+ 513,    8*2048+ 958,    0*2048+1141,
  18*2048+  36,   34*2048+ 992,   44*2048+1014,    0*2048+1142,
  28*2048+ 120,   38*2048+ 306,   11*2048+ 613,    0*2048+1147,
  38*2048+ 609,   12*2048+ 680,   20*2048+ 898,    0*2048+1148,
  43*2048+ 263,   42*2048+ 624,    5*2048+ 645,    0*2048+1149,
   9*2048+  13,   22*2048+ 394,   15*2048+ 649,    0*2048+1150,
  35*2048+  48,   45*2048+  69,   18*2048+ 171,    0*2048+1151,
  22*2048+  43,    1*2048+  60,   17*2048+ 151,   19*2048+ 357,   33*2048+ 459,    0*2048+ 540,   43*2048+ 648,   26*2048+ 777,    5*2048+ 826,   16*2048+ 867,   21*2048+ 925,   38*2048+ 972,    0*2048+1080,
  28*2048+  20,   37*2048+ 131,   12*2048+ 143,   17*2048+ 346,   13*2048+ 432,   38*2048+ 548,   10*2048+ 718,   26*2048+ 747,   20*2048+ 766,   28*2048+ 870,   35*2048+ 874,   12*2048+1044,    0*2048+1081,
  18*2048+  91,   25*2048+ 147,    9*2048+ 309,   12*2048+ 349,   30*2048+ 397,   37*2048+ 444,   12*2048+ 591,   42*2048+ 635,   26*2048+ 706,   38*2048+ 875,   22*2048+ 926,   14*2048+ 976,    0*2048+1082,
  17*2048+  47,    9*2048+ 132,   41*2048+ 230,   32*2048+ 258,   30*2048+ 294,   36*2048+ 350,   11*2048+ 623,   38*2048+ 659,   23*2048+ 679,   20*2048+ 830,   12*2048+ 945,   36*2048+1057,    0*2048+1083,
  39*2048+  27,   22*2048+ 178,    1*2048+ 195,   17*2048+ 286,   19*2048+ 492,   33*2048+ 594,    0*2048+ 675,   43*2048+ 784,   26*2048+ 912,    5*2048+ 961,   16*2048+1002,   21*2048+1060,    0*2048+1089,
  13*2048+  99,   28*2048+ 155,   37*2048+ 266,   12*2048+ 278,   17*2048+ 481,   13*2048+ 567,   38*2048+ 683,   10*2048+ 853,   26*2048+ 882,   20*2048+ 901,   28*2048+1005,   35*2048+1009,    0*2048+1090,
  15*2048+  31,   18*2048+ 226,   25*2048+ 282,    9*2048+ 445,   12*2048+ 484,   30*2048+ 532,   37*2048+ 579,   12*2048+ 726,   42*2048+ 770,   26*2048+ 841,   38*2048+1010,   22*2048+1061,    0*2048+1091,
  13*2048+   0,   37*2048+ 112,   17*2048+ 183,    9*2048+ 267,   41*2048+ 365,   32*2048+ 393,   30*2048+ 429,   36*2048+ 485,   11*2048+ 759,   38*2048+ 794,   23*2048+ 815,   20*2048+ 965,    0*2048+1092,
   6*2048+  16,   17*2048+  57,   22*2048+ 115,   39*2048+ 162,   22*2048+ 313,    1*2048+ 330,   17*2048+ 421,   19*2048+ 627,   33*2048+ 729,    0*2048+ 810,   43*2048+ 919,   26*2048+1047,    0*2048+1098,
  29*2048+  61,   36*2048+  64,   13*2048+ 234,   28*2048+ 290,   37*2048+ 401,   12*2048+ 413,   17*2048+ 616,   13*2048+ 702,   38*2048+ 818,   10*2048+ 988,   26*2048+1017,   20*2048+1036,    0*2048+1099,
  39*2048+  65,   23*2048+ 116,   15*2048+ 166,   18*2048+ 361,   25*2048+ 417,    9*2048+ 580,   12*2048+ 619,   30*2048+ 667,   37*2048+ 714,   12*2048+ 861,   42*2048+ 905,   26*2048+ 977,    0*2048+1100,
  21*2048+  21,   13*2048+ 135,   37*2048+ 247,   17*2048+ 318,    9*2048+ 402,   41*2048+ 500,   32*2048+ 529,   30*2048+ 564,   36*2048+ 620,   11*2048+ 894,   38*2048+ 929,   23*2048+ 950,    0*2048+1101,
  27*2048+ 102,    6*2048+ 152,   17*2048+ 192,   22*2048+ 250,   39*2048+ 297,   22*2048+ 448,    1*2048+ 465,   17*2048+ 556,   19*2048+ 762,   33*2048+ 864,    0*2048+ 946,   43*2048+1054,    0*2048+1107,
  11*2048+  44,   27*2048+  72,   21*2048+  92,   29*2048+ 196,   36*2048+ 199,   13*2048+ 369,   28*2048+ 425,   37*2048+ 536,   12*2048+ 549,   17*2048+ 751,   13*2048+ 837,   38*2048+ 953,    0*2048+1108,
  27*2048+  32,   39*2048+ 200,   23*2048+ 251,   15*2048+ 301,   18*2048+ 496,   25*2048+ 552,    9*2048+ 715,   12*2048+ 754,   30*2048+ 802,   37*2048+ 849,   12*2048+ 996,   42*2048+1040,    0*2048+1109,
  24*2048+   5,   21*2048+ 156,   13*2048+ 270,   37*2048+ 382,   17*2048+ 453,    9*2048+ 537,   41*2048+ 636,   32*2048+ 664,   30*2048+ 699,   36*2048+ 755,   11*2048+1029,   38*2048+1064,    0*2048+1110,
   1*2048+   1,   44*2048+ 109,   27*2048+ 237,    6*2048+ 287,   17*2048+ 327,   22*2048+ 385,   39*2048+ 433,   22*2048+ 583,    1*2048+ 600,   17*2048+ 691,   19*2048+ 897,   33*2048+ 999,    0*2048+1116,
  39*2048+   8,   11*2048+ 179,   27*2048+ 207,   21*2048+ 227,   29*2048+ 331,   36*2048+ 334,   13*2048+ 504,   28*2048+ 560,   37*2048+ 671,   12*2048+ 684,   17*2048+ 886,   13*2048+ 973,    0*2048+1117,
  13*2048+  51,   43*2048+  95,   27*2048+ 167,   39*2048+ 335,   23*2048+ 386,   15*2048+ 436,   18*2048+ 631,   25*2048+ 687,    9*2048+ 850,   12*2048+ 889,   30*2048+ 937,   37*2048+ 984,    0*2048+1118,
  12*2048+  84,   39*2048+ 119,   24*2048+ 140,   21*2048+ 291,   13*2048+ 405,   37*2048+ 517,   17*2048+ 588,    9*2048+ 672,   41*2048+ 771,   32*2048+ 799,   30*2048+ 834,   36*2048+ 890,    0*2048+1119,
  34*2048+  54,    1*2048+ 136,   44*2048+ 244,   27*2048+ 372,    6*2048+ 422,   17*2048+ 462,   22*2048+ 520,   39*2048+ 568,   22*2048+ 719,    1*2048+ 735,   17*2048+ 827,   19*2048+1033,    0*2048+1125,
  14*2048+  28,   39*2048+ 144,   11*2048+ 314,   27*2048+ 342,   21*2048+ 362,   29*2048+ 466,   36*2048+ 469,   13*2048+ 639,   28*2048+ 695,   37*2048+ 806,   12*2048+ 819,   17*2048+1021,    0*2048+1126,
  38*2048+  39,   13*2048+ 186,   43*2048+ 231,   27*2048+ 302,   39*2048+ 470,   23*2048+ 521,   15*2048+ 571,   18*2048+ 767,   25*2048+ 822,    9*2048+ 985,   12*2048+1024,   30*2048+1072,    0*2048+1127,
  12*2048+ 219,   39*2048+ 255,   24*2048+ 275,   21*2048+ 426,   13*2048+ 541,   37*2048+ 652,   17*2048+ 723,    9*2048+ 807,   41*2048+ 906,   32*2048+ 934,   30*2048+ 969,   36*2048+1025,    0*2048+1128,
  20*2048+  88,   34*2048+ 189,    1*2048+ 271,   44*2048+ 379,   27*2048+ 507,    6*2048+ 557,   17*2048+ 597,   22*2048+ 655,   39*2048+ 703,   22*2048+ 854,    1*2048+ 871,   17*2048+ 962,    0*2048+1134,
  18*2048+  76,   14*2048+ 163,   39*2048+ 279,   11*2048+ 449,   27*2048+ 477,   21*2048+ 497,   29*2048+ 601,   36*2048+ 604,   13*2048+ 774,   28*2048+ 831,   37*2048+ 941,   12*2048+ 954,    0*2048+1135,
  10*2048+  40,   13*2048+  79,   31*2048+ 127,   38*2048+ 174,   13*2048+ 321,   43*2048+ 366,   27*2048+ 437,   39*2048+ 605,   23*2048+ 656,   15*2048+ 707,   18*2048+ 902,   25*2048+ 957,    0*2048+1136,
  31*2048+  24,   37*2048+  80,   12*2048+ 354,   39*2048+ 390,   24*2048+ 410,   21*2048+ 561,   13*2048+ 676,   37*2048+ 787,   17*2048+ 858,    9*2048+ 942,   41*2048+1041,   32*2048+1069,    0*2048+1137,
  18*2048+  17,   20*2048+ 223,   34*2048+ 324,    1*2048+ 406,   44*2048+ 514,   27*2048+ 642,    6*2048+ 692,   17*2048+ 732,   22*2048+ 790,   39*2048+ 838,   22*2048+ 989,    1*2048+1006,    0*2048+1143,
  13*2048+   9,   18*2048+ 211,   14*2048+ 298,   39*2048+ 414,   11*2048+ 584,   27*2048+ 612,   21*2048+ 632,   29*2048+ 736,   36*2048+ 739,   13*2048+ 909,   28*2048+ 966,   37*2048+1076,    0*2048+1144,
  26*2048+  12,   10*2048+ 175,   13*2048+ 214,   31*2048+ 262,   38*2048+ 310,   13*2048+ 456,   43*2048+ 501,   27*2048+ 572,   39*2048+ 740,   23*2048+ 791,   15*2048+ 842,   18*2048+1037,    0*2048+1145,
  42*2048+  96,   33*2048+ 124,   31*2048+ 159,   37*2048+ 215,   12*2048+ 489,   39*2048+ 525,   24*2048+ 545,   21*2048+ 696,   13*2048+ 811,   37*2048+ 922,   17*2048+ 993,    9*2048+1077,    0*2048+1146,

   0*2048+   3,    0*2048+   8,    0*2048+1320,
   0*2048+   9,    0*2048+  13,    0*2048+1321,
   0*2048+  14,    0*2048+  18,    0*2048+1322,
   0*2048+  19,    0*2048+  23,    0*2048+1323,
   0*2048+  24,    0*2048+  28,    0*2048+1324,
   0*2048+  29,    0*2048+  33,    0*2048+1325,
   0*2048+  34,    0*2048+  38,    0*2048+1326,
   0*2048+  39,    0*2048+  43,    0*2048+1327,
   0*2048+  44,    0*2048+  48,    0*2048+1328,
   0*2048+  49,    0*2048+  53,    0*2048+1329,
   0*2048+  54,    0*2048+  58,    0*2048+1330,
   0*2048+  59,    0*2048+  63,    0*2048+1331,
   0*2048+  64,    0*2048+  68,    0*2048+1332,
   0*2048+  69,    0*2048+  73,    0*2048+1333,
   0*2048+  74,    0*2048+  78,    0*2048+1334,
   0*2048+  79,    0*2048+  83,    0*2048+1335,
   0*2048+  84,    0*2048+  88,    0*2048+1336,
   0*2048+  89,    0*2048+  93,    0*2048+1337,
   0*2048+  94,    0*2048+  98,    0*2048+1338,
   0*2048+  99,    0*2048+ 103,    0*2048+1339,
   0*2048+ 104,    0*2048+ 108,    0*2048+1340,
   0*2048+ 109,    0*2048+ 113,    0*2048+1341,
   0*2048+ 114,    0*2048+ 118,    0*2048+1342,
   0*2048+ 119,    0*2048+ 123,    0*2048+1343,
   0*2048+ 124,    0*2048+ 128,    0*2048+1344,
   0*2048+ 129,    0*2048+ 133,    0*2048+1345,
   0*2048+ 134,    0*2048+ 138,    0*2048+1346,
   0*2048+ 139,    0*2048+ 143,    0*2048+1347,
   0*2048+ 144,    0*2048+ 148,    0*2048+1348,
   0*2048+ 149,    0*2048+ 153,    0*2048+1349,
   0*2048+ 154,    0*2048+ 158,    0*2048+1350,
   0*2048+ 159,    0*2048+ 163,    0*2048+1351,
   0*2048+ 164,    0*2048+ 168,    0*2048+1352,
   0*2048+ 169,    0*2048+ 173,    0*2048+1353,
   0*2048+ 174,    0*2048+ 178,    0*2048+1354,
   0*2048+ 179,    0*2048+ 183,    0*2048+1355,
   0*2048+ 184,    0*2048+ 188,    0*2048+1356,
   0*2048+ 189,    0*2048+ 193,    0*2048+1357,
   0*2048+ 194,    0*2048+ 198,    0*2048+1358,
   0*2048+ 199,    0*2048+ 203,    0*2048+1359,
   0*2048+ 204,    0*2048+ 208,    0*2048+1360,
   0*2048+ 209,    0*2048+ 213,    0*2048+1361,
   0*2048+ 214,    0*2048+ 218,    0*2048+1362,
   0*2048+ 219,    0*2048+ 223,    0*2048+1363,
   0*2048+ 224,    0*2048+ 228,    0*2048+1364,
   0*2048+ 229,    0*2048+ 233,    0*2048+1365,
   0*2048+ 234,    0*2048+ 238,    0*2048+1366,
   0*2048+ 239,    0*2048+ 243,    0*2048+1367,
   0*2048+ 244,    0*2048+ 248,    0*2048+1368,
   0*2048+ 249,    0*2048+ 253,    0*2048+1369,
   0*2048+ 254,    0*2048+ 258,    0*2048+1370,
   0*2048+ 259,    0*2048+ 263,    0*2048+1371,
   0*2048+ 264,    0*2048+ 268,    0*2048+1372,
   0*2048+ 269,    0*2048+ 273,    0*2048+1373,
   0*2048+ 274,    0*2048+ 278,    0*2048+1374,
   0*2048+ 279,    0*2048+ 283,    0*2048+1375,
   0*2048+ 284,    0*2048+ 288,    0*2048+1376,
   0*2048+ 289,    0*2048+ 293,    0*2048+1377,
   0*2048+ 294,    0*2048+ 298,    0*2048+1378,
   0*2048+ 299,    0*2048+ 303,    0*2048+1379,
   0*2048+ 304,    0*2048+ 308,    0*2048+1380,
   0*2048+ 309,    0*2048+ 313,    0*2048+1381,
   0*2048+ 314,    0*2048+ 318,    0*2048+1382,
   0*2048+ 319,    0*2048+ 323,    0*2048+1383,
   0*2048+ 324,    0*2048+ 328,    0*2048+1384,
   0*2048+ 329,    0*2048+ 333,    0*2048+1385,
   0*2048+ 334,    0*2048+ 338,    0*2048+1386,
   0*2048+ 339,    0*2048+ 343,    0*2048+1387,
   0*2048+ 344,    0*2048+ 348,    0*2048+1388,
   0*2048+ 349,    0*2048+ 353,    0*2048+1389,
   0*2048+ 354,    0*2048+ 358,    0*2048+1390,
   0*2048+ 359,    0*2048+ 363,    0*2048+1391,
   0*2048+ 364,    0*2048+ 368,    0*2048+1392,
   0*2048+ 369,    0*2048+ 373,    0*2048+1393,
   0*2048+ 374,    0*2048+ 378,    0*2048+1394,
   0*2048+ 379,    0*2048+ 383,    0*2048+1395,
   0*2048+ 384,    0*2048+ 388,    0*2048+1396,
   0*2048+ 389,    0*2048+ 393,    0*2048+1397,
   0*2048+ 394,    0*2048+ 398,    0*2048+1398,
   0*2048+ 399,    0*2048+ 403,    0*2048+1399,
   0*2048+ 404,    0*2048+ 408,    0*2048+1400,
   0*2048+ 409,    0*2048+ 413,    0*2048+1401,
   0*2048+ 414,    0*2048+ 418,    0*2048+1402,
   0*2048+ 419,    0*2048+ 423,    0*2048+1403,
   0*2048+ 424,    0*2048+ 428,    0*2048+1404,
   0*2048+ 429,    0*2048+ 433,    0*2048+1405,
   0*2048+ 434,    0*2048+ 438,    0*2048+1406,
   0*2048+ 439,    0*2048+ 443,    0*2048+1407,
   0*2048+ 444,    0*2048+ 448,    0*2048+1408,
   0*2048+ 449,    0*2048+ 453,    0*2048+1409,
   0*2048+ 454,    0*2048+ 458,    0*2048+1410,
   0*2048+ 459,    0*2048+ 463,    0*2048+1411,
   0*2048+ 464,    0*2048+ 468,    0*2048+1412,
   0*2048+ 469,    0*2048+ 473,    0*2048+1413,
   0*2048+ 474,    0*2048+ 478,    0*2048+1414,
   0*2048+ 479,    0*2048+ 483,    0*2048+1415,
   0*2048+ 484,    0*2048+ 488,    0*2048+1416,
   0*2048+ 489,    0*2048+ 493,    0*2048+1417,
   0*2048+ 494,    0*2048+ 498,    0*2048+1418,
   0*2048+ 499,    0*2048+ 503,    0*2048+1419,
   0*2048+ 504,    0*2048+ 508,    0*2048+1420,
   0*2048+ 509,    0*2048+ 513,    0*2048+1421,
   0*2048+ 514,    0*2048+ 518,    0*2048+1422,
   0*2048+ 519,    0*2048+ 523,    0*2048+1423,
   0*2048+ 524,    0*2048+ 528,    0*2048+1424,
   0*2048+ 529,    0*2048+ 533,    0*2048+1425,
   0*2048+ 534,    0*2048+ 538,    0*2048+1426,
   0*2048+ 539,    0*2048+ 543,    0*2048+1427,
   0*2048+ 544,    0*2048+ 548,    0*2048+1428,
   0*2048+ 549,    0*2048+ 553,    0*2048+1429,
   0*2048+ 554,    0*2048+ 558,    0*2048+1430,
   0*2048+ 559,    0*2048+ 563,    0*2048+1431,
   0*2048+ 564,    0*2048+ 568,    0*2048+1432,
   0*2048+ 569,    0*2048+ 573,    0*2048+1433,
   0*2048+ 574,    0*2048+ 578,    0*2048+1434,
   0*2048+ 579,    0*2048+ 583,    0*2048+1435,
   0*2048+ 584,    0*2048+ 588,    0*2048+1436,
   0*2048+ 589,    0*2048+ 593,    0*2048+1437,
   0*2048+ 594,    0*2048+ 598,    0*2048+1438,
   0*2048+ 599,    0*2048+ 603,    0*2048+1439,
   0*2048+ 604,    0*2048+ 608,    0*2048+1440,
   0*2048+ 609,    0*2048+ 613,    0*2048+1441,
   0*2048+ 614,    0*2048+ 618,    0*2048+1442,
   0*2048+ 619,    0*2048+ 623,    0*2048+1443,
   0*2048+ 624,    0*2048+ 628,    0*2048+1444,
   0*2048+ 629,    0*2048+ 633,    0*2048+1445,
   0*2048+ 634,    0*2048+ 638,    0*2048+1446,
   0*2048+ 639,    0*2048+ 643,    0*2048+1447,
   0*2048+ 644,    0*2048+ 648,    0*2048+1448,
   0*2048+ 649,    0*2048+ 653,    0*2048+1449,
   0*2048+ 654,    0*2048+ 658,    0*2048+1450,
   0*2048+ 659,    0*2048+ 663,    0*2048+1451,
   0*2048+ 664,    0*2048+ 668,    0*2048+1452,
   0*2048+ 669,    0*2048+ 673,    0*2048+1453,
   0*2048+ 674,    0*2048+ 678,    0*2048+1454,
   0*2048+ 679,    0*2048+ 683,    0*2048+1455,
   0*2048+ 684,    0*2048+ 688,    0*2048+1456,
   0*2048+ 689,    0*2048+ 693,    0*2048+1457,
   0*2048+ 694,    0*2048+ 698,    0*2048+1458,
   0*2048+ 699,    0*2048+ 703,    0*2048+1459,
   0*2048+ 704,    0*2048+ 708,    0*2048+1460,
   0*2048+ 709,    0*2048+ 713,    0*2048+1461,
   0*2048+ 714,    0*2048+ 718,    0*2048+1462,
   0*2048+ 719,    0*2048+ 723,    0*2048+1463,
   0*2048+ 724,    0*2048+ 728,    0*2048+1464,
   0*2048+ 729,    0*2048+ 733,    0*2048+1465,
   0*2048+ 734,    0*2048+ 738,    0*2048+1466,
   0*2048+ 739,    0*2048+ 743,    0*2048+1467,
   0*2048+ 744,    0*2048+ 748,    0*2048+1468,
   0*2048+ 749,    0*2048+ 753,    0*2048+1469,
   0*2048+ 754,    0*2048+ 758,    0*2048+1470,
   0*2048+ 759,    0*2048+ 763,    0*2048+1471,
   0*2048+ 764,    0*2048+ 768,    0*2048+1472,
   0*2048+ 769,    0*2048+ 773,    0*2048+1473,
   0*2048+ 774,    0*2048+ 778,    0*2048+1474,
   0*2048+ 779,    0*2048+ 783,    0*2048+1475,
   0*2048+ 784,    0*2048+ 788,    0*2048+1476,
   0*2048+ 789,    0*2048+ 793,    0*2048+1477,
   0*2048+ 794,    0*2048+ 798,    0*2048+1478,
   0*2048+ 799,    0*2048+ 803,    0*2048+1479,
   0*2048+ 804,    0*2048+ 808,    0*2048+1480,
   0*2048+ 809,    0*2048+ 813,    0*2048+1481,
   0*2048+ 814,    0*2048+ 818,    0*2048+1482,
   0*2048+ 819,    0*2048+ 823,    0*2048+1483,
   0*2048+ 824,    0*2048+ 828,    0*2048+1484,
   0*2048+ 829,    0*2048+ 833,    0*2048+1485,
   0*2048+ 834,    0*2048+ 838,    0*2048+1486,
   0*2048+ 839,    0*2048+ 843,    0*2048+1487,
   0*2048+ 844,    0*2048+ 848,    0*2048+1488,
   0*2048+ 849,    0*2048+ 853,    0*2048+1489,
   0*2048+ 854,    0*2048+ 858,    0*2048+1490,
   0*2048+ 859,    0*2048+ 863,    0*2048+1491,
   0*2048+ 864,    0*2048+ 868,    0*2048+1492,
   0*2048+ 869,    0*2048+ 873,    0*2048+1493,
   0*2048+ 874,    0*2048+ 878,    0*2048+1494,
   0*2048+ 879,    0*2048+ 883,    0*2048+1495,
   0*2048+ 884,    0*2048+ 888,    0*2048+1496,
   0*2048+ 889,    0*2048+ 893,    0*2048+1497,
   0*2048+ 894,    0*2048+ 898,    0*2048+1498,
   0*2048+ 899,    0*2048+ 903,    0*2048+1499,
   0*2048+ 904,    0*2048+ 908,    0*2048+1500,
   0*2048+ 909,    0*2048+ 913,    0*2048+1501,
   0*2048+ 914,    0*2048+ 918,    0*2048+1502,
   0*2048+ 919,    0*2048+ 923,    0*2048+1503,
   0*2048+ 924,    0*2048+ 928,    0*2048+1504,
   0*2048+ 929,    0*2048+ 933,    0*2048+1505,
   0*2048+ 934,    0*2048+ 938,    0*2048+1506,
   0*2048+ 939,    0*2048+ 943,    0*2048+1507,
   0*2048+ 944,    0*2048+ 948,    0*2048+1508,
   0*2048+ 949,    0*2048+ 953,    0*2048+1509,
   0*2048+ 954,    0*2048+ 958,    0*2048+1510,
   0*2048+ 959,    0*2048+ 963,    0*2048+1511,
   0*2048+ 964,    0*2048+ 968,    0*2048+1512,
   0*2048+ 969,    0*2048+ 973,    0*2048+1513,
   0*2048+ 974,    0*2048+ 978,    0*2048+1514,
   0*2048+ 979,    0*2048+ 983,    0*2048+1515,
   0*2048+ 984,    0*2048+ 988,    0*2048+1516,
   0*2048+ 989,    0*2048+ 993,    0*2048+1517,
   0*2048+ 994,    0*2048+ 998,    0*2048+1518,
   0*2048+ 999,    0*2048+1003,    0*2048+1519,
   0*2048+1004,    0*2048+1008,    0*2048+1520,
   0*2048+1009,    0*2048+1013,    0*2048+1521,
   0*2048+1014,    0*2048+1018,    0*2048+1522,
   0*2048+1019,    0*2048+1023,    0*2048+1523,
   0*2048+1024,    0*2048+1028,    0*2048+1524,
   0*2048+1029,    0*2048+1033,    0*2048+1525,
   0*2048+1034,    0*2048+1038,    0*2048+1526,
   0*2048+1039,    0*2048+1043,    0*2048+1527,
   0*2048+1044,    0*2048+1048,    0*2048+1528,
   0*2048+1049,    0*2048+1053,    0*2048+1529,
   0*2048+1054,    0*2048+1058,    0*2048+1530,
   0*2048+1059,    0*2048+1063,    0*2048+1531,
   0*2048+1064,    0*2048+1068,    0*2048+1532,
   0*2048+1069,    0*2048+1073,    0*2048+1533,
   0*2048+1074,    0*2048+1078,    0*2048+1534,
   0*2048+1079,    0*2048+1083,    0*2048+1535,
   0*2048+1084,    0*2048+1088,    0*2048+1536,
   0*2048+1089,    0*2048+1093,    0*2048+1537,
   0*2048+1094,    0*2048+1098,    0*2048+1538,
   0*2048+1099,    0*2048+1103,    0*2048+1539,
   0*2048+1104,    0*2048+1108,    0*2048+1540,
   0*2048+1109,    0*2048+1113,    0*2048+1541,
   0*2048+1114,    0*2048+1118,    0*2048+1542,
   0*2048+1119,    0*2048+1123,    0*2048+1543,
   0*2048+1124,    0*2048+1128,    0*2048+1544,
   0*2048+1129,    0*2048+1133,    0*2048+1545,
   0*2048+1134,    0*2048+1138,    0*2048+1546,
   0*2048+1139,    0*2048+1143,    0*2048+1547,
   0*2048+1144,    0*2048+1148,    0*2048+1548,
   0*2048+1149,    0*2048+1153,    0*2048+1549,
   0*2048+1154,    0*2048+1158,    0*2048+1550,
   0*2048+1159,    0*2048+1163,    0*2048+1551,
   0*2048+1164,    0*2048+1168,    0*2048+1552,
   0*2048+1169,    0*2048+1173,    0*2048+1553,
   0*2048+1174,    0*2048+1178,    0*2048+1554,
   0*2048+1179,    0*2048+1183,    0*2048+1555,
   0*2048+1184,    0*2048+1188,    0*2048+1556,
   0*2048+1189,    0*2048+1193,    0*2048+1557,
   0*2048+1194,    0*2048+1198,    0*2048+1558,
   1*2048+   4,    0*2048+1199,    0*2048+1559,
   6*2048+ 325,   32*2048+ 491,   23*2048+ 810,    0*2048+1205,
  28*2048+ 551,   27*2048+ 715,   29*2048+1060,    0*2048+1206,
  30*2048+ 406,   16*2048+ 505,   14*2048+ 725,    0*2048+1207,
  36*2048+ 146,   42*2048+ 950,    3*2048+ 971,    0*2048+1208,
  15*2048+ 111,   39*2048+ 140,   31*2048+ 615,    0*2048+1209,
  21*2048+  90,   41*2048+ 450,   18*2048+1170,    0*2048+1210,
  40*2048+  45,   20*2048+ 220,   11*2048+ 336,    0*2048+1211,
   7*2048+ 170,   13*2048+ 586,   28*2048+ 815,    0*2048+1212,
  16*2048+ 190,   41*2048+ 885,   19*2048+1040,    0*2048+1213,
  42*2048+ 235,   34*2048+ 535,   13*2048+1070,    0*2048+1214,
   6*2048+ 475,   32*2048+ 641,   23*2048+ 962,    0*2048+1220,
  30*2048+  10,   28*2048+ 702,   27*2048+ 865,    0*2048+1221,
  30*2048+ 556,   16*2048+ 657,   14*2048+ 876,    0*2048+1222,
  36*2048+ 296,   42*2048+1100,    3*2048+1121,    0*2048+1223,
  15*2048+ 261,   39*2048+ 290,   31*2048+ 765,    0*2048+1224,
  19*2048+ 121,   21*2048+ 240,   41*2048+ 600,    0*2048+1225,
  40*2048+ 195,   20*2048+ 370,   11*2048+ 486,    0*2048+1226,
   7*2048+ 320,   13*2048+ 736,   28*2048+ 966,    0*2048+1227,
  16*2048+ 340,   41*2048+1035,   19*2048+1190,    0*2048+1228,
  14*2048+  20,   42*2048+ 386,   34*2048+ 685,    0*2048+1229,
   6*2048+ 625,   32*2048+ 791,   23*2048+1112,    0*2048+1235,
  30*2048+ 161,   28*2048+ 852,   27*2048+1015,    0*2048+1236,
  30*2048+ 706,   16*2048+ 807,   14*2048+1027,    0*2048+1237,
  43*2048+  50,    4*2048+  71,   36*2048+ 446,    0*2048+1238,
  15*2048+ 411,   39*2048+ 441,   31*2048+ 915,    0*2048+1239,
  19*2048+ 271,   21*2048+ 390,   41*2048+ 750,    0*2048+1240,
  40*2048+ 345,   20*2048+ 520,   11*2048+ 636,    0*2048+1241,
   7*2048+ 470,   13*2048+ 887,   28*2048+1116,    0*2048+1242,
  20*2048+ 141,   16*2048+ 492,   41*2048+1185,    0*2048+1243,
  14*2048+ 171,   42*2048+ 537,   34*2048+ 835,    0*2048+1244,
  24*2048+  62,    6*2048+ 775,   32*2048+ 941,    0*2048+1250,
  30*2048+ 311,   28*2048+1002,   27*2048+1165,    0*2048+1251,
  30*2048+ 856,   16*2048+ 957,   14*2048+1177,    0*2048+1252,
  43*2048+ 200,    4*2048+ 222,   36*2048+ 596,    0*2048+1253,
  15*2048+ 561,   39*2048+ 591,   31*2048+1065,    0*2048+1254,
  19*2048+ 421,   21*2048+ 540,   41*2048+ 900,    0*2048+1255,
  40*2048+ 496,   20*2048+ 670,   11*2048+ 787,    0*2048+1256,
  29*2048+  66,    7*2048+ 620,   13*2048+1037,    0*2048+1257,
  42*2048+ 135,   20*2048+ 291,   16*2048+ 642,    0*2048+1258,
  14*2048+ 321,   42*2048+ 687,   34*2048+ 985,    0*2048+1259,
  24*2048+ 212,    6*2048+ 925,   32*2048+1091,    0*2048+1265,
  28*2048+ 117,   30*2048+ 461,   28*2048+1152,    0*2048+1266,
  15*2048+ 127,   30*2048+1006,   16*2048+1107,    0*2048+1267,
  43*2048+ 350,    4*2048+ 372,   36*2048+ 746,    0*2048+1268,
  32*2048+  16,   15*2048+ 711,   39*2048+ 741,    0*2048+1269,
  19*2048+ 571,   21*2048+ 691,   41*2048+1051,    0*2048+1270,
  40*2048+ 646,   20*2048+ 820,   11*2048+ 937,    0*2048+1271,
  29*2048+ 216,    7*2048+ 771,   13*2048+1187,    0*2048+1272,
  42*2048+ 285,   20*2048+ 442,   16*2048+ 792,    0*2048+1273,
  14*2048+ 471,   42*2048+ 837,   34*2048+1135,    0*2048+1274,
  33*2048+  41,   24*2048+ 362,    6*2048+1077,    0*2048+1280,
  29*2048+ 102,   28*2048+ 267,   30*2048+ 611,    0*2048+1281,
  17*2048+  57,   15*2048+ 277,   30*2048+1156,    0*2048+1282,
  43*2048+ 501,    4*2048+ 522,   36*2048+ 896,    0*2048+1283,
  32*2048+ 166,   15*2048+ 861,   39*2048+ 891,    0*2048+1284,
  42*2048+   2,   19*2048+ 721,   21*2048+ 842,    0*2048+1285,
  40*2048+ 796,   20*2048+ 972,   11*2048+1087,    0*2048+1286,
  14*2048+ 137,   29*2048+ 366,    7*2048+ 921,    0*2048+1287,
  42*2048+ 435,   20*2048+ 592,   16*2048+ 942,    0*2048+1288,
  35*2048+  85,   14*2048+ 621,   42*2048+ 987,    0*2048+1289,
   7*2048+  27,   33*2048+ 192,   24*2048+ 512,    0*2048+1295,
  29*2048+ 252,   28*2048+ 417,   30*2048+ 762,    0*2048+1296,
  31*2048+ 107,   17*2048+ 207,   15*2048+ 427,    0*2048+1297,
  43*2048+ 651,    4*2048+ 672,   36*2048+1047,    0*2048+1298,
  32*2048+ 316,   15*2048+1011,   39*2048+1042,    0*2048+1299,
  42*2048+ 152,   19*2048+ 871,   21*2048+ 992,    0*2048+1300,
  12*2048+  37,   40*2048+ 946,   20*2048+1122,    0*2048+1301,
  14*2048+ 287,   29*2048+ 517,    7*2048+1072,    0*2048+1302,
  42*2048+ 587,   20*2048+ 742,   16*2048+1092,    0*2048+1303,
  35*2048+ 236,   14*2048+ 772,   42*2048+1137,    0*2048+1304,
   7*2048+ 177,   33*2048+ 342,   24*2048+ 662,    0*2048+1310,
  29*2048+ 402,   28*2048+ 567,   30*2048+ 912,    0*2048+1311,
  31*2048+ 257,   17*2048+ 357,   15*2048+ 577,    0*2048+1312,
  43*2048+ 802,    4*2048+ 822,   36*2048+1197,    0*2048+1313,
  32*2048+ 467,   15*2048+1162,   39*2048+1192,    0*2048+1314,
  42*2048+ 302,   19*2048+1022,   21*2048+1142,    0*2048+1315,
  21*2048+  72,   12*2048+ 187,   40*2048+1097,    0*2048+1316,
   8*2048+  22,   14*2048+ 437,   29*2048+ 667,    0*2048+1317,
  17*2048+  42,   42*2048+ 737,   20*2048+ 892,    0*2048+1318,
  43*2048+  87,   35*2048+ 387,   14*2048+ 922,    0*2048+1319,
  28*2048+  15,   37*2048+ 145,   12*2048+ 160,   17*2048+ 380,   13*2048+ 480,   10*2048+ 800,   26*2048+ 825,   20*2048+ 845,    1*2048+ 880,   28*2048+ 960,   35*2048+ 965,   12*2048+1160,    0*2048+1200,
  18*2048+  95,   25*2048+ 155,    9*2048+ 330,   12*2048+ 385,   30*2048+ 440,   37*2048+ 490,   12*2048+ 655,   42*2048+ 690,   26*2048+ 780,   38*2048+ 961,   22*2048+1025,   14*2048+1075,    0*2048+1201,
  14*2048+ 115,   39*2048+ 120,    8*2048+ 225,   42*2048+ 335,   21*2048+ 495,    9*2048+ 656,    4*2048+ 770,   41*2048+ 840,   14*2048+ 881,    1*2048+ 970,   17*2048+1050,   41*2048+1095,    0*2048+1202,
  16*2048+   0,    8*2048+ 105,   19*2048+ 110,    3*2048+ 116,   36*2048+ 381,   15*2048+ 465,   21*2048+ 500,   29*2048+ 585,   22*2048+ 700,   11*2048+ 785,   31*2048+ 875,   25*2048+1076,    0*2048+1203,
   6*2048+ 375,   20*2048+ 395,   14*2048+ 405,   22*2048+ 515,   25*2048+ 550,   20*2048+ 730,   35*2048+ 755,    7*2048+ 756,   43*2048+ 760,   30*2048+1020,   39*2048+1045,   17*2048+1130,    0*2048+1204,
  13*2048+ 112,   28*2048+ 165,   37*2048+ 295,   12*2048+ 310,   17*2048+ 530,   13*2048+ 630,   10*2048+ 951,   26*2048+ 975,   20*2048+ 995,    1*2048+1030,   28*2048+1110,   35*2048+1115,    0*2048+1215,
  15*2048+  25,   18*2048+ 245,   25*2048+ 305,    9*2048+ 481,   12*2048+ 536,   30*2048+ 590,   37*2048+ 640,   12*2048+ 805,   42*2048+ 841,   26*2048+ 930,   38*2048+1111,   22*2048+1175,    0*2048+1216,
  18*2048+   1,   42*2048+  46,   14*2048+ 265,   39*2048+ 270,    8*2048+ 376,   42*2048+ 485,   21*2048+ 645,    9*2048+ 806,    4*2048+ 920,   41*2048+ 990,   14*2048+1031,    1*2048+1120,    0*2048+1217,
  26*2048+  26,   16*2048+ 150,    8*2048+ 255,   19*2048+ 260,    3*2048+ 266,   36*2048+ 531,   15*2048+ 616,   21*2048+ 650,   29*2048+ 735,   22*2048+ 850,   11*2048+ 935,   31*2048+1026,    0*2048+1218,
  18*2048+  80,    6*2048+ 525,   20*2048+ 545,   14*2048+ 555,   22*2048+ 665,   25*2048+ 701,   20*2048+ 882,   35*2048+ 905,    7*2048+ 906,   43*2048+ 910,   30*2048+1171,   39*2048+1195,    0*2048+1219,
  29*2048+  60,   36*2048+  65,   13*2048+ 262,   28*2048+ 315,   37*2048+ 445,   12*2048+ 460,   17*2048+ 680,   13*2048+ 781,   10*2048+1101,   26*2048+1125,   20*2048+1145,    1*2048+1180,    0*2048+1230,
  39*2048+  61,   23*2048+ 125,   15*2048+ 175,   18*2048+ 396,   25*2048+ 455,    9*2048+ 631,   12*2048+ 686,   30*2048+ 740,   37*2048+ 790,   12*2048+ 955,   42*2048+ 991,   26*2048+1080,    0*2048+1231,
   2*2048+  70,   18*2048+ 151,   42*2048+ 196,   14*2048+ 415,   39*2048+ 420,    8*2048+ 526,   42*2048+ 635,   21*2048+ 795,    9*2048+ 956,    4*2048+1071,   41*2048+1140,   14*2048+1181,    0*2048+1232,
  26*2048+ 176,   16*2048+ 300,    8*2048+ 407,   19*2048+ 410,    3*2048+ 416,   36*2048+ 681,   15*2048+ 766,   21*2048+ 801,   29*2048+ 886,   22*2048+1000,   11*2048+1085,   31*2048+1176,    0*2048+1233,
  31*2048+ 122,   40*2048+ 147,   18*2048+ 230,    6*2048+ 675,   20*2048+ 695,   14*2048+ 705,   22*2048+ 816,   25*2048+ 851,   20*2048+1032,   35*2048+1055,    7*2048+1056,   43*2048+1061,    0*2048+1234,
  11*2048+  51,   27*2048+  75,   21*2048+  96,    2*2048+ 130,   29*2048+ 210,   36*2048+ 215,   13*2048+ 412,   28*2048+ 466,   37*2048+ 595,   12*2048+ 610,   17*2048+ 830,   13*2048+ 931,    0*2048+1245,
  27*2048+  30,   39*2048+ 211,   23*2048+ 275,   15*2048+ 326,   18*2048+ 546,   25*2048+ 605,    9*2048+ 782,   12*2048+ 836,   30*2048+ 890,   37*2048+ 940,   12*2048+1105,   42*2048+1141,    0*2048+1246,
   5*2048+  21,   42*2048+  91,   15*2048+ 131,    2*2048+ 221,   18*2048+ 301,   42*2048+ 346,   14*2048+ 565,   39*2048+ 570,    8*2048+ 676,   42*2048+ 786,   21*2048+ 945,    9*2048+1106,    0*2048+1247,
  12*2048+  35,   32*2048+ 126,   26*2048+ 327,   16*2048+ 451,    8*2048+ 557,   19*2048+ 560,    3*2048+ 566,   36*2048+ 831,   15*2048+ 916,   21*2048+ 952,   29*2048+1036,   22*2048+1150,    0*2048+1248,
  36*2048+   5,    8*2048+   6,   44*2048+  11,   31*2048+ 272,   40*2048+ 297,   18*2048+ 382,    6*2048+ 826,   20*2048+ 846,   14*2048+ 855,   22*2048+ 967,   25*2048+1001,   20*2048+1182,    0*2048+1249,
  11*2048+ 201,   27*2048+ 226,   21*2048+ 246,    2*2048+ 280,   29*2048+ 360,   36*2048+ 365,   13*2048+ 562,   28*2048+ 617,   37*2048+ 745,   12*2048+ 761,   17*2048+ 980,   13*2048+1081,    0*2048+1260,
  13*2048+  55,   43*2048+  92,   27*2048+ 180,   39*2048+ 361,   23*2048+ 425,   15*2048+ 476,   18*2048+ 696,   25*2048+ 757,    9*2048+ 932,   12*2048+ 986,   30*2048+1041,   37*2048+1090,    0*2048+1261,
  10*2048+  56,    5*2048+ 172,   42*2048+ 241,   15*2048+ 281,    2*2048+ 371,   18*2048+ 452,   42*2048+ 497,   14*2048+ 716,   39*2048+ 720,    8*2048+ 827,   42*2048+ 936,   21*2048+1096,    0*2048+1262,
  23*2048+ 100,   12*2048+ 185,   32*2048+ 276,   26*2048+ 477,   16*2048+ 601,    8*2048+ 707,   19*2048+ 710,    3*2048+ 717,   36*2048+ 981,   15*2048+1066,   21*2048+1102,   29*2048+1186,    0*2048+1263,
  21*2048+ 132,   36*2048+ 156,    8*2048+ 157,   44*2048+ 162,   31*2048+ 422,   40*2048+ 447,   18*2048+ 532,    6*2048+ 976,   20*2048+ 996,   14*2048+1005,   22*2048+1117,   25*2048+1151,    0*2048+1264,
  14*2048+  31,   11*2048+ 351,   27*2048+ 377,   21*2048+ 397,    2*2048+ 430,   29*2048+ 510,   36*2048+ 516,   13*2048+ 712,   28*2048+ 767,   37*2048+ 895,   12*2048+ 911,   17*2048+1131,    0*2048+1275,
  38*2048+  40,   13*2048+ 205,   43*2048+ 242,   27*2048+ 331,   39*2048+ 511,   23*2048+ 575,   15*2048+ 626,   18*2048+ 847,   25*2048+ 907,    9*2048+1082,   12*2048+1136,   30*2048+1191,    0*2048+1276,
  22*2048+  47,   10*2048+ 206,    5*2048+ 322,   42*2048+ 391,   15*2048+ 431,    2*2048+ 521,   18*2048+ 602,   42*2048+ 647,   14*2048+ 866,   39*2048+ 870,    8*2048+ 977,   42*2048+1086,    0*2048+1277,
  16*2048+  17,   22*2048+  52,   30*2048+ 136,   23*2048+ 250,   12*2048+ 337,   32*2048+ 426,   26*2048+ 627,   16*2048+ 751,    8*2048+ 857,   19*2048+ 860,    3*2048+ 867,   36*2048+1132,    0*2048+1278,
  23*2048+  67,   26*2048+ 101,   21*2048+ 282,   36*2048+ 306,    8*2048+ 307,   44*2048+ 312,   31*2048+ 572,   40*2048+ 597,   18*2048+ 682,    6*2048+1126,   20*2048+1146,   14*2048+1155,    0*2048+1279,
  18*2048+  81,   14*2048+ 181,   11*2048+ 502,   27*2048+ 527,   21*2048+ 547,    2*2048+ 580,   29*2048+ 660,   36*2048+ 666,   13*2048+ 862,   28*2048+ 917,   37*2048+1046,   12*2048+1062,    0*2048+1290,
  10*2048+  32,   13*2048+  86,   31*2048+ 142,   38*2048+ 191,   13*2048+ 355,   43*2048+ 392,   27*2048+ 482,   39*2048+ 661,   23*2048+ 726,   15*2048+ 776,   18*2048+ 997,   25*2048+1057,    0*2048+1291,
  43*2048+  36,   22*2048+ 197,   10*2048+ 356,    5*2048+ 472,   42*2048+ 541,   15*2048+ 581,    2*2048+ 671,   18*2048+ 752,   42*2048+ 797,   14*2048+1016,   39*2048+1021,    8*2048+1127,    0*2048+1292,
  37*2048+  82,   16*2048+ 167,   22*2048+ 202,   30*2048+ 286,   23*2048+ 400,   12*2048+ 487,   32*2048+ 576,   26*2048+ 777,   16*2048+ 901,    8*2048+1007,   19*2048+1010,    3*2048+1017,    0*2048+1293,
   7*2048+  76,   21*2048+  97,   15*2048+ 106,   23*2048+ 217,   26*2048+ 251,   21*2048+ 432,   36*2048+ 456,    8*2048+ 457,   44*2048+ 462,   31*2048+ 722,   40*2048+ 747,   18*2048+ 832,    0*2048+1294,
  13*2048+  12,   18*2048+ 231,   14*2048+ 332,   11*2048+ 652,   27*2048+ 677,   21*2048+ 697,    2*2048+ 731,   29*2048+ 811,   36*2048+ 817,   13*2048+1012,   28*2048+1067,   37*2048+1196,    0*2048+1305,
  26*2048+   7,   10*2048+ 182,   13*2048+ 237,   31*2048+ 292,   38*2048+ 341,   13*2048+ 506,   43*2048+ 542,   27*2048+ 632,   39*2048+ 812,   23*2048+ 877,   15*2048+ 926,   18*2048+1147,    0*2048+1306,
   9*2048+  77,   43*2048+ 186,   22*2048+ 347,   10*2048+ 507,    5*2048+ 622,   42*2048+ 692,   15*2048+ 732,    2*2048+ 821,   18*2048+ 902,   42*2048+ 947,   14*2048+1166,   39*2048+1172,    0*2048+1307,
  37*2048+ 232,   16*2048+ 317,   22*2048+ 352,   30*2048+ 436,   23*2048+ 552,   12*2048+ 637,   32*2048+ 727,   26*2048+ 927,   16*2048+1052,    8*2048+1157,   19*2048+1161,    3*2048+1167,    0*2048+1308,
   7*2048+ 227,   21*2048+ 247,   15*2048+ 256,   23*2048+ 367,   26*2048+ 401,   21*2048+ 582,   36*2048+ 606,    8*2048+ 607,   44*2048+ 612,   31*2048+ 872,   40*2048+ 897,   18*2048+ 982,    0*2048+1309,

   0*2048+   4,    0*2048+  10,    0*2048+1440,
   0*2048+  11,    0*2048+  16,    0*2048+1441,
   0*2048+  17,    0*2048+  22,    0*2048+1442,
   0*2048+  23,    0*2048+  28,    0*2048+1443,
   0*2048+  29,    0*2048+  34,    0*2048+1444,
   0*2048+  35,    0*2048+  40,    0*2048+1445,
   0*2048+  41,    0*2048+  46,    0*2048+1446,
   0*2048+  47,    0*2048+  52,    0*2048+1447,
   0*2048+  53,    0*2048+  58,    0*2048+1448,
   0*2048+  59,    0*2048+  64,    0*2048+1449,
   0*2048+  65,    0*2048+  70,    0*2048+1450,
   0*2048+  71,    0*2048+  76,    0*2048+1451,
   0*2048+  77,    0*2048+  82,    0*2048+1452,
   0*2048+  83,    0*2048+  88,    0*2048+1453,
   0*2048+  89,    0*2048+  94,    0*2048+1454,
   0*2048+  95,    0*2048+ 100,    0*2048+1455,
   0*2048+ 101,    0*2048+ 106,    0*2048+1456,
   0*2048+ 107,    0*2048+ 112,    0*2048+1457,
   0*2048+ 113,    0*2048+ 118,    0*2048+1458,
   0*2048+ 119,    0*2048+ 124,    0*2048+1459,
   0*2048+ 125,    0*2048+ 130,    0*2048+1460,
   0*2048+ 131,    0*2048+ 136,    0*2048+1461,
   0*2048+ 137,    0*2048+ 142,    0*2048+1462,
   0*2048+ 143,    0*2048+ 148,    0*2048+1463,
   0*2048+ 149,    0*2048+ 154,    0*2048+1464,
   0*2048+ 155,    0*2048+ 160,    0*2048+1465,
   0*2048+ 161,    0*2048+ 166,    0*2048+1466,
   0*2048+ 167,    0*2048+ 172,    0*2048+1467,
   0*2048+ 173,    0*2048+ 178,    0*2048+1468,
   0*2048+ 179,    0*2048+ 184,    0*2048+1469,
   0*2048+ 185,    0*2048+ 190,    0*2048+1470,
   0*2048+ 191,    0*2048+ 196,    0*2048+1471,
   0*2048+ 197,    0*2048+ 202,    0*2048+1472,
   0*2048+ 203,    0*2048+ 208,    0*2048+1473,
   0*2048+ 209,    0*2048+ 214,    0*2048+1474,
   0*2048+ 215,    0*2048+ 220,    0*2048+1475,
   0*2048+ 221,    0*2048+ 226,    0*2048+1476,
   0*2048+ 227,    0*2048+ 232,    0*2048+1477,
   0*2048+ 233,    0*2048+ 238,    0*2048+1478,
   0*2048+ 239,    0*2048+ 244,    0*2048+1479,
   0*2048+ 245,    0*2048+ 250,    0*2048+1480,
   0*2048+ 251,    0*2048+ 256,    0*2048+1481,
   0*2048+ 257,    0*2048+ 262,    0*2048+1482,
   0*2048+ 263,    0*2048+ 268,    0*2048+1483,
   0*2048+ 269,    0*2048+ 274,    0*2048+1484,
   0*2048+ 275,    0*2048+ 280,    0*2048+1485,
   0*2048+ 281,    0*2048+ 286,    0*2048+1486,
   0*2048+ 287,    0*2048+ 292,    0*2048+1487,
   0*2048+ 293,    0*2048+ 298,    0*2048+1488,
   0*2048+ 299,    0*2048+ 304,    0*2048+1489,
   0*2048+ 305,    0*2048+ 310,    0*2048+1490,
   0*2048+ 311,    0*2048+ 316,    0*2048+1491,
   0*2048+ 317,    0*2048+ 322,    0*2048+1492,
   0*2048+ 323,    0*2048+ 328,    0*2048+1493,
   0*2048+ 329,    0*2048+ 334,    0*2048+1494,
   0*2048+ 335,    0*2048+ 340,    0*2048+1495,
   0*2048+ 341,    0*2048+ 346,    0*2048+1496,
   0*2048+ 347,    0*2048+ 352,    0*2048+1497,
   0*2048+ 353,    0*2048+ 358,    0*2048+1498,
   0*2048+ 359,    0*2048+ 364,    0*2048+1499,
   0*2048+ 365,    0*2048+ 370,    0*2048+1500,
   0*2048+ 371,    0*2048+ 376,    0*2048+1501,
   0*2048+ 377,    0*2048+ 382,    0*2048+1502,
   0*2048+ 383,    0*2048+ 388,    0*2048+1503,
   0*2048+ 389,    0*2048+ 394,    0*2048+1504,
   0*2048+ 395,    0*2048+ 400,    0*2048+1505,
   0*2048+ 401,    0*2048+ 406,    0*2048+1506,
   0*2048+ 407,    0*2048+ 412,    0*2048+1507,
   0*2048+ 413,    0*2048+ 418,    0*2048+1508,
   0*2048+ 419,    0*2048+ 424,    0*2048+1509,
   0*2048+ 425,    0*2048+ 430,    0*2048+1510,
   0*2048+ 431,    0*2048+ 436,    0*2048+1511,
   0*2048+ 437,    0*2048+ 442,    0*2048+1512,
   0*2048+ 443,    0*2048+ 448,    0*2048+1513,
   0*2048+ 449,    0*2048+ 454,    0*2048+1514,
   0*2048+ 455,    0*2048+ 460,    0*2048+1515,
   0*2048+ 461,    0*2048+ 466,    0*2048+1516,
   0*2048+ 467,    0*2048+ 472,    0*2048+1517,
   0*2048+ 473,    0*2048+ 478,    0*2048+1518,
   0*2048+ 479,    0*2048+ 484,    0*2048+1519,
   0*2048+ 485,    0*2048+ 490,    0*2048+1520,
   0*2048+ 491,    0*2048+ 496,    0*2048+1521,
   0*2048+ 497,    0*2048+ 502,    0*2048+1522,
   0*2048+ 503,    0*2048+ 508,    0*2048+1523,
   0*2048+ 509,    0*2048+ 514,    0*2048+1524,
   0*2048+ 515,    0*2048+ 520,    0*2048+1525,
   0*2048+ 521,    0*2048+ 526,    0*2048+1526,
   0*2048+ 527,    0*2048+ 532,    0*2048+1527,
   0*2048+ 533,    0*2048+ 538,    0*2048+1528,
   0*2048+ 539,    0*2048+ 544,    0*2048+1529,
   0*2048+ 545,    0*2048+ 550,    0*2048+1530,
   0*2048+ 551,    0*2048+ 556,    0*2048+1531,
   0*2048+ 557,    0*2048+ 562,    0*2048+1532,
   0*2048+ 563,    0*2048+ 568,    0*2048+1533,
   0*2048+ 569,    0*2048+ 574,    0*2048+1534,
   0*2048+ 575,    0*2048+ 580,    0*2048+1535,
   0*2048+ 581,    0*2048+ 586,    0*2048+1536,
   0*2048+ 587,    0*2048+ 592,    0*2048+1537,
   0*2048+ 593,    0*2048+ 598,    0*2048+1538,
   0*2048+ 599,    0*2048+ 604,    0*2048+1539,
   0*2048+ 605,    0*2048+ 610,    0*2048+1540,
   0*2048+ 611,    0*2048+ 616,    0*2048+1541,
   0*2048+ 617,    0*2048+ 622,    0*2048+1542,
   0*2048+ 623,    0*2048+ 628,    0*2048+1543,
   0*2048+ 629,    0*2048+ 634,    0*2048+1544,
   0*2048+ 635,    0*2048+ 640,    0*2048+1545,
   0*2048+ 641,    0*2048+ 646,    0*2048+1546,
   0*2048+ 647,    0*2048+ 652,    0*2048+1547,
   0*2048+ 653,    0*2048+ 658,    0*2048+1548,
   0*2048+ 659,    0*2048+ 664,    0*2048+1549,
   0*2048+ 665,    0*2048+ 670,    0*2048+1550,
   0*2048+ 671,    0*2048+ 676,    0*2048+1551,
   0*2048+ 677,    0*2048+ 682,    0*2048+1552,
   0*2048+ 683,    0*2048+ 688,    0*2048+1553,
   0*2048+ 689,    0*2048+ 694,    0*2048+1554,
   0*2048+ 695,    0*2048+ 700,    0*2048+1555,
   0*2048+ 701,    0*2048+ 706,    0*2048+1556,
   0*2048+ 707,    0*2048+ 712,    0*2048+1557,
   0*2048+ 713,    0*2048+ 718,    0*2048+1558,
   0*2048+ 719,    0*2048+ 724,    0*2048+1559,
   0*2048+ 725,    0*2048+ 730,    0*2048+1560,
   0*2048+ 731,    0*2048+ 736,    0*2048+1561,
   0*2048+ 737,    0*2048+ 742,    0*2048+1562,
   0*2048+ 743,    0*2048+ 748,    0*2048+1563,
   0*2048+ 749,    0*2048+ 754,    0*2048+1564,
   0*2048+ 755,    0*2048+ 760,    0*2048+1565,
   0*2048+ 761,    0*2048+ 766,    0*2048+1566,
   0*2048+ 767,    0*2048+ 772,    0*2048+1567,
   0*2048+ 773,    0*2048+ 778,    0*2048+1568,
   0*2048+ 779,    0*2048+ 784,    0*2048+1569,
   0*2048+ 785,    0*2048+ 790,    0*2048+1570,
   0*2048+ 791,    0*2048+ 796,    0*2048+1571,
   0*2048+ 797,    0*2048+ 802,    0*2048+1572,
   0*2048+ 803,    0*2048+ 808,    0*2048+1573,
   0*2048+ 809,    0*2048+ 814,    0*2048+1574,
   0*2048+ 815,    0*2048+ 820,    0*2048+1575,
   0*2048+ 821,    0*2048+ 826,    0*2048+1576,
   0*2048+ 827,    0*2048+ 832,    0*2048+1577,
   0*2048+ 833,    0*2048+ 838,    0*2048+1578,
   0*2048+ 839,    0*2048+ 844,    0*2048+1579,
   0*2048+ 845,    0*2048+ 850,    0*2048+1580,
   0*2048+ 851,    0*2048+ 856,    0*2048+1581,
   0*2048+ 857,    0*2048+ 862,    0*2048+1582,
   0*2048+ 863,    0*2048+ 868,    0*2048+1583,
   0*2048+ 869,    0*2048+ 874,    0*2048+1584,
   0*2048+ 875,    0*2048+ 880,    0*2048+1585,
   0*2048+ 881,    0*2048+ 886,    0*2048+1586,
   0*2048+ 887,    0*2048+ 892,    0*2048+1587,
   0*2048+ 893,    0*2048+ 898,    0*2048+1588,
   0*2048+ 899,    0*2048+ 904,    0*2048+1589,
   0*2048+ 905,    0*2048+ 910,    0*2048+1590,
   0*2048+ 911,    0*2048+ 916,    0*2048+1591,
   0*2048+ 917,    0*2048+ 922,    0*2048+1592,
   0*2048+ 923,    0*2048+ 928,    0*2048+1593,
   0*2048+ 929,    0*2048+ 934,    0*2048+1594,
   0*2048+ 935,    0*2048+ 940,    0*2048+1595,
   0*2048+ 941,    0*2048+ 946,    0*2048+1596,
   0*2048+ 947,    0*2048+ 952,    0*2048+1597,
   0*2048+ 953,    0*2048+ 958,    0*2048+1598,
   0*2048+ 959,    0*2048+ 964,    0*2048+1599,
   0*2048+ 965,    0*2048+ 970,    0*2048+1600,
   0*2048+ 971,    0*2048+ 976,    0*2048+1601,
   0*2048+ 977,    0*2048+ 982,    0*2048+1602,
   0*2048+ 983,    0*2048+ 988,    0*2048+1603,
   0*2048+ 989,    0*2048+ 994,    0*2048+1604,
   0*2048+ 995,    0*2048+1000,    0*2048+1605,
   0*2048+1001,    0*2048+1006,    0*2048+1606,
   0*2048+1007,    0*2048+1012,    0*2048+1607,
   0*2048+1013,    0*2048+1018,    0*2048+1608,
   0*2048+1019,    0*2048+1024,    0*2048+1609,
   0*2048+1025,    0*2048+1030,    0*2048+1610,
   0*2048+1031,    0*2048+1036,    0*2048+1611,
   0*2048+1037,    0*2048+1042,    0*2048+1612,
   0*2048+1043,    0*2048+1048,    0*2048+1613,
   0*2048+1049,    0*2048+1054,    0*2048+1614,
   0*2048+1055,    0*2048+1060,    0*2048+1615,
   0*2048+1061,    0*2048+1066,    0*2048+1616,
   0*2048+1067,    0*2048+1072,    0*2048+1617,
   0*2048+1073,    0*2048+1078,    0*2048+1618,
   0*2048+1079,    0*2048+1084,    0*2048+1619,
   0*2048+1085,    0*2048+1090,    0*2048+1620,
   0*2048+1091,    0*2048+1096,    0*2048+1621,
   0*2048+1097,    0*2048+1102,    0*2048+1622,
   0*2048+1103,    0*2048+1108,    0*2048+1623,
   0*2048+1109,    0*2048+1114,    0*2048+1624,
   0*2048+1115,    0*2048+1120,    0*2048+1625,
   0*2048+1121,    0*2048+1126,    0*2048+1626,
   0*2048+1127,    0*2048+1132,    0*2048+1627,
   0*2048+1133,    0*2048+1138,    0*2048+1628,
   0*2048+1139,    0*2048+1144,    0*2048+1629,
   0*2048+1145,    0*2048+1150,    0*2048+1630,
   0*2048+1151,    0*2048+1156,    0*2048+1631,
   0*2048+1157,    0*2048+1162,    0*2048+1632,
   0*2048+1163,    0*2048+1168,    0*2048+1633,
   0*2048+1169,    0*2048+1174,    0*2048+1634,
   0*2048+1175,    0*2048+1180,    0*2048+1635,
   0*2048+1181,    0*2048+1186,    0*2048+1636,
   0*2048+1187,    0*2048+1192,    0*2048+1637,
   0*2048+1193,    0*2048+1198,    0*2048+1638,
   0*2048+1199,    0*2048+1204,    0*2048+1639,
   0*2048+1205,    0*2048+1210,    0*2048+1640,
   0*2048+1211,    0*2048+1216,    0*2048+1641,
   0*2048+1217,    0*2048+1222,    0*2048+1642,
   0*2048+1223,    0*2048+1228,    0*2048+1643,
   0*2048+1229,    0*2048+1234,    0*2048+1644,
   0*2048+1235,    0*2048+1240,    0*2048+1645,
   0*2048+1241,    0*2048+1246,    0*2048+1646,
   0*2048+1247,    0*2048+1252,    0*2048+1647,
   0*2048+1253,    0*2048+1258,    0*2048+1648,
   0*2048+1259,    0*2048+1264,    0*2048+1649,
   0*2048+1265,    0*2048+1270,    0*2048+1650,
   0*2048+1271,    0*2048+1276,    0*2048+1651,
   0*2048+1277,    0*2048+1282,    0*2048+1652,
   0*2048+1283,    0*2048+1288,    0*2048+1653,
   0*2048+1289,    0*2048+1294,    0*2048+1654,
   1*2048+   5,    0*2048+1295,    0*2048+1655,
   6*2048+ 834,    7*2048+ 840,   37*2048+1074,    0*2048+1302,
  30*2048+ 378,   17*2048+ 438,   15*2048+ 756,    0*2048+1303,
  39*2048+ 510,   21*2048+ 655,   42*2048+1284,    0*2048+1304,
  34*2048+ 318,   41*2048+ 696,   26*2048+1044,    0*2048+1305,
   8*2048+ 426,   20*2048+ 612,   30*2048+ 702,    0*2048+1306,
  18*2048+ 918,   17*2048+1050,   42*2048+1224,    0*2048+1307,
  34*2048+ 206,   40*2048+ 258,   22*2048+1164,    0*2048+1308,
   9*2048+ 294,   42*2048+ 686,   24*2048+ 984,    0*2048+1309,
  31*2048+ 168,   26*2048+ 181,   41*2048+ 954,    0*2048+1310,
  39*2048+ 300,   20*2048+ 714,   20*2048+1092,    0*2048+1311,
  23*2048+ 835,   43*2048+ 924,   33*2048+1285,    0*2048+1312,
  41*2048+ 324,   12*2048+ 409,    6*2048+ 546,    0*2048+1313,
   6*2048+ 996,    7*2048+1002,   37*2048+1237,    0*2048+1320,
  30*2048+ 541,   17*2048+ 600,   15*2048+ 919,    0*2048+1321,
  43*2048+ 150,   39*2048+ 672,   21*2048+ 817,    0*2048+1322,
  34*2048+ 481,   41*2048+ 859,   26*2048+1207,    0*2048+1323,
   8*2048+ 588,   20*2048+ 774,   30*2048+ 865,    0*2048+1324,
  43*2048+  90,   18*2048+1080,   17*2048+1212,    0*2048+1325,
  23*2048+  30,   34*2048+ 368,   40*2048+ 420,    0*2048+1326,
   9*2048+ 456,   42*2048+ 849,   24*2048+1146,    0*2048+1327,
  31*2048+ 331,   26*2048+ 343,   41*2048+1116,    0*2048+1328,
  39*2048+ 462,   20*2048+ 876,   20*2048+1255,    0*2048+1329,
  34*2048+ 151,   23*2048+ 997,   43*2048+1087,    0*2048+1330,
  41*2048+ 486,   12*2048+ 571,    6*2048+ 708,    0*2048+1331,
  38*2048+ 104,    6*2048+1158,    7*2048+1165,    0*2048+1338,
  30*2048+ 704,   17*2048+ 762,   15*2048+1081,    0*2048+1339,
  43*2048+ 312,   39*2048+ 836,   21*2048+ 979,    0*2048+1340,
  27*2048+  73,   34*2048+ 645,   41*2048+1021,    0*2048+1341,
   8*2048+ 750,   20*2048+ 937,   30*2048+1027,    0*2048+1342,
  18*2048+  79,   43*2048+ 254,   18*2048+1242,    0*2048+1343,
  23*2048+ 193,   34*2048+ 530,   40*2048+ 582,    0*2048+1344,
  25*2048+  12,    9*2048+ 618,   42*2048+1011,    0*2048+1345,
  31*2048+ 493,   26*2048+ 505,   41*2048+1278,    0*2048+1346,
  21*2048+ 121,   39*2048+ 625,   20*2048+1039,    0*2048+1347,
  34*2048+ 313,   23*2048+1159,   43*2048+1250,    0*2048+1348,
  41*2048+ 650,   12*2048+ 733,    6*2048+ 870,    0*2048+1349,
   7*2048+  25,    8*2048+  31,   38*2048+ 266,    0*2048+1356,
  30*2048+ 867,   17*2048+ 925,   15*2048+1243,    0*2048+1357,
  43*2048+ 475,   39*2048+ 998,   21*2048+1141,    0*2048+1358,
  27*2048+ 237,   34*2048+ 807,   41*2048+1183,    0*2048+1359,
   8*2048+ 912,   20*2048+1100,   30*2048+1189,    0*2048+1360,
  19*2048+ 109,   18*2048+ 241,   43*2048+ 416,    0*2048+1361,
  23*2048+ 355,   34*2048+ 692,   40*2048+ 744,    0*2048+1362,
  25*2048+ 174,    9*2048+ 781,   42*2048+1173,    0*2048+1363,
  42*2048+ 147,   31*2048+ 657,   26*2048+ 667,    0*2048+1364,
  21*2048+ 284,   39*2048+ 787,   20*2048+1202,    0*2048+1365,
  24*2048+  26,   44*2048+ 116,   34*2048+ 476,    0*2048+1366,
  41*2048+ 812,   12*2048+ 895,    6*2048+1033,    0*2048+1367,
   7*2048+ 187,    8*2048+ 194,   38*2048+ 429,    0*2048+1374,
  16*2048+ 110,   30*2048+1029,   17*2048+1088,    0*2048+1375,
  22*2048+   7,   43*2048+ 637,   39*2048+1160,    0*2048+1376,
  42*2048+  49,   27*2048+ 399,   34*2048+ 969,    0*2048+1377,
  31*2048+  55,    8*2048+1075,   20*2048+1262,    0*2048+1378,
  19*2048+ 271,   18*2048+ 404,   43*2048+ 578,    0*2048+1379,
  23*2048+ 517,   34*2048+ 855,   40*2048+ 907,    0*2048+1380,
  43*2048+  39,   25*2048+ 336,    9*2048+ 943,    0*2048+1381,
  42*2048+ 309,   31*2048+ 819,   26*2048+ 830,    0*2048+1382,
  21*2048+  69,   21*2048+ 447,   39*2048+ 950,    0*2048+1383,
  24*2048+ 188,   44*2048+ 278,   34*2048+ 638,    0*2048+1384,
  41*2048+ 974,   12*2048+1057,    6*2048+1196,    0*2048+1385,
   7*2048+ 349,    8*2048+ 356,   38*2048+ 591,    0*2048+1392,
  16*2048+ 272,   30*2048+1191,   17*2048+1251,    0*2048+1393,
  40*2048+  27,   22*2048+ 170,   43*2048+ 799,    0*2048+1394,
  42*2048+ 212,   27*2048+ 561,   34*2048+1131,    0*2048+1395,
  21*2048+ 128,   31*2048+ 217,    8*2048+1238,    0*2048+1396,
  19*2048+ 434,   18*2048+ 567,   43*2048+ 741,    0*2048+1397,
  23*2048+ 680,   34*2048+1017,   40*2048+1070,    0*2048+1398,
  43*2048+ 201,   25*2048+ 499,    9*2048+1105,    0*2048+1399,
  42*2048+ 471,   31*2048+ 981,   26*2048+ 992,    0*2048+1400,
  21*2048+ 231,   21*2048+ 609,   39*2048+1112,    0*2048+1401,
  24*2048+ 350,   44*2048+ 441,   34*2048+ 800,    0*2048+1402,
   7*2048+  63,   41*2048+1137,   12*2048+1221,    0*2048+1403,
   7*2048+ 512,    8*2048+ 518,   38*2048+ 753,    0*2048+1410,
  31*2048+  57,   18*2048+ 117,   16*2048+ 435,    0*2048+1411,
  40*2048+ 189,   22*2048+ 333,   43*2048+ 961,    0*2048+1412,
  42*2048+ 374,   27*2048+ 723,   34*2048+1293,    0*2048+1413,
   9*2048+ 105,   21*2048+ 291,   31*2048+ 380,    0*2048+1414,
  19*2048+ 596,   18*2048+ 729,   43*2048+ 903,    0*2048+1415,
  23*2048+ 843,   34*2048+1179,   40*2048+1232,    0*2048+1416,
  43*2048+ 363,   25*2048+ 663,    9*2048+1267,    0*2048+1417,
  42*2048+ 633,   31*2048+1143,   26*2048+1154,    0*2048+1418,
  21*2048+ 393,   21*2048+ 771,   39*2048+1275,    0*2048+1419,
  24*2048+ 513,   44*2048+ 603,   34*2048+ 962,    0*2048+1420,
  42*2048+   3,   13*2048+  87,    7*2048+ 225,    0*2048+1421,
   7*2048+ 674,    8*2048+ 681,   38*2048+ 915,    0*2048+1428,
  31*2048+ 219,   18*2048+ 279,   16*2048+ 597,    0*2048+1429,
  40*2048+ 351,   22*2048+ 495,   43*2048+1124,    0*2048+1430,
  35*2048+ 159,   42*2048+ 537,   27*2048+ 885,    0*2048+1431,
   9*2048+ 267,   21*2048+ 453,   31*2048+ 543,    0*2048+1432,
  19*2048+ 759,   18*2048+ 891,   43*2048+1065,    0*2048+1433,
  35*2048+  45,   41*2048+  99,   23*2048+1005,    0*2048+1434,
  10*2048+ 135,   43*2048+ 525,   25*2048+ 825,    0*2048+1435,
  32*2048+   9,   27*2048+  21,   42*2048+ 795,    0*2048+1436,
  40*2048+ 141,   21*2048+ 555,   21*2048+ 933,    0*2048+1437,
  24*2048+ 675,   44*2048+ 765,   34*2048+1125,    0*2048+1438,
  42*2048+ 165,   13*2048+ 249,    7*2048+ 387,    0*2048+1439,
  32*2048+  60,   31*2048+ 144,   26*2048+ 204,   19*2048+ 234,    8*2048+ 235,    6*2048+ 288,   37*2048+ 474,    3*2048+ 540,   40*2048+ 660,    2*2048+ 906,   30*2048+1068,    2*2048+1218,    0*2048+1296,
  32*2048+  18,   12*2048+  78,   37*2048+ 145,    8*2048+ 252,   23*2048+ 330,   26*2048+ 480,   32*2048+ 642,    7*2048+1038,   14*2048+1098,    1*2048+1194,   25*2048+1248,    3*2048+1254,    0*2048+1297,
  36*2048+  96,    4*2048+ 132,   10*2048+ 180,    8*2048+ 444,   28*2048+ 534,   18*2048+ 624,   41*2048+ 684,    3*2048+ 738,   33*2048+ 780,    8*2048+ 828,   40*2048+1206,    8*2048+1219,    0*2048+1298,
  19*2048+  24,   35*2048+ 102,   38*2048+ 108,   43*2048+ 205,   27*2048+ 210,   10*2048+ 564,   20*2048+ 648,   17*2048+ 654,   31*2048+ 685,   40*2048+1122,   35*2048+1236,   24*2048+1272,    0*2048+1299,
   1*2048+  66,   22*2048+ 133,    4*2048+ 146,   27*2048+ 192,   20*2048+ 282,   41*2048+ 643,    1*2048+ 649,   36*2048+ 678,   29*2048+ 846,   19*2048+ 858,   44*2048+ 936,   40*2048+1086,    0*2048+1300,
  43*2048+ 253,   10*2048+ 402,    2*2048+ 408,   22*2048+ 432,    8*2048+ 498,   14*2048+ 661,   18*2048+ 852,   11*2048+ 864,    3*2048+ 948,   23*2048+1032,   44*2048+1134,    8*2048+1200,    0*2048+1301,
   3*2048+  84,   32*2048+ 222,   31*2048+ 306,   26*2048+ 366,   19*2048+ 396,    8*2048+ 397,    6*2048+ 450,   37*2048+ 636,    3*2048+ 703,   40*2048+ 822,    2*2048+1069,   30*2048+1230,    0*2048+1314,
   2*2048+  61,   26*2048+ 114,    4*2048+ 120,   32*2048+ 182,   12*2048+ 240,   37*2048+ 307,    8*2048+ 414,   23*2048+ 492,   26*2048+ 644,   32*2048+ 804,    7*2048+1201,   14*2048+1260,    0*2048+1315,
  41*2048+  72,    9*2048+  85,   36*2048+ 259,    4*2048+ 295,   10*2048+ 342,    8*2048+ 606,   28*2048+ 697,   18*2048+ 786,   41*2048+ 847,    3*2048+ 900,   33*2048+ 942,    8*2048+ 990,    0*2048+1316,
  36*2048+ 103,   25*2048+ 138,   19*2048+ 186,   35*2048+ 264,   38*2048+ 270,   43*2048+ 367,   27*2048+ 372,   10*2048+ 726,   20*2048+ 810,   17*2048+ 816,   31*2048+ 848,   40*2048+1286,    0*2048+1317,
   1*2048+ 228,   22*2048+ 296,    4*2048+ 308,   27*2048+ 354,   20*2048+ 445,   41*2048+ 805,    1*2048+ 811,   36*2048+ 841,   29*2048+1008,   19*2048+1020,   44*2048+1099,   40*2048+1249,    0*2048+1318,
  45*2048+   0,    9*2048+  67,   43*2048+ 415,   10*2048+ 565,    2*2048+ 570,   22*2048+ 594,    8*2048+ 662,   14*2048+ 823,   18*2048+1014,   11*2048+1026,    3*2048+1110,   23*2048+1195,    0*2048+1319,
  31*2048+  97,    3*2048+ 246,   32*2048+ 384,   31*2048+ 468,   26*2048+ 528,   19*2048+ 558,    8*2048+ 559,    6*2048+ 613,   37*2048+ 798,    3*2048+ 866,   40*2048+ 985,    2*2048+1231,    0*2048+1332,
   8*2048+  68,   15*2048+ 126,    2*2048+ 223,   26*2048+ 276,    4*2048+ 283,   32*2048+ 344,   12*2048+ 403,   37*2048+ 469,    8*2048+ 576,   23*2048+ 656,   26*2048+ 806,   32*2048+ 966,    0*2048+1333,
  41*2048+ 236,    9*2048+ 247,   36*2048+ 421,    4*2048+ 457,   10*2048+ 504,    8*2048+ 768,   28*2048+ 860,   18*2048+ 949,   41*2048+1009,    3*2048+1062,   33*2048+1104,    8*2048+1152,    0*2048+1334,
  41*2048+ 152,   36*2048+ 265,   25*2048+ 301,   19*2048+ 348,   35*2048+ 427,   38*2048+ 433,   43*2048+ 529,   27*2048+ 535,   10*2048+ 888,   20*2048+ 972,   17*2048+ 978,   31*2048+1010,    0*2048+1335,
  41*2048+ 115,    1*2048+ 390,   22*2048+ 458,    4*2048+ 470,   27*2048+ 516,   20*2048+ 607,   41*2048+ 967,    1*2048+ 973,   36*2048+1003,   29*2048+1170,   19*2048+1182,   44*2048+1261,    0*2048+1336,
  24*2048+  62,   45*2048+ 162,    9*2048+ 229,   43*2048+ 577,   10*2048+ 727,    2*2048+ 732,   22*2048+ 757,    8*2048+ 824,   14*2048+ 986,   18*2048+1176,   11*2048+1188,    3*2048+1273,    0*2048+1337,
   3*2048+  98,   31*2048+ 260,    3*2048+ 410,   32*2048+ 547,   31*2048+ 630,   26*2048+ 690,   19*2048+ 720,    8*2048+ 721,    6*2048+ 775,   37*2048+ 960,    3*2048+1028,   40*2048+1147,    0*2048+1350,
   8*2048+ 230,   15*2048+ 289,    2*2048+ 385,   26*2048+ 439,    4*2048+ 446,   32*2048+ 506,   12*2048+ 566,   37*2048+ 631,    8*2048+ 739,   23*2048+ 818,   26*2048+ 968,   32*2048+1128,    0*2048+1351,
   9*2048+  19,   41*2048+ 398,    9*2048+ 411,   36*2048+ 583,    4*2048+ 619,   10*2048+ 666,    8*2048+ 930,   28*2048+1022,   18*2048+1111,   41*2048+1171,    3*2048+1225,   33*2048+1266,    0*2048+1352,
  41*2048+ 314,   36*2048+ 428,   25*2048+ 463,   19*2048+ 511,   35*2048+ 589,   38*2048+ 595,   43*2048+ 691,   27*2048+ 698,   10*2048+1051,   20*2048+1135,   17*2048+1140,   31*2048+1172,    0*2048+1353,
  30*2048+  36,   20*2048+  48,   45*2048+ 127,   41*2048+ 277,    1*2048+ 552,   22*2048+ 620,    4*2048+ 632,   27*2048+ 679,   20*2048+ 769,   41*2048+1129,    1*2048+1136,   36*2048+1166,    0*2048+1354,
  19*2048+  42,   12*2048+  54,    4*2048+ 139,   24*2048+ 224,   45*2048+ 325,    9*2048+ 391,   43*2048+ 740,   10*2048+ 889,    2*2048+ 894,   22*2048+ 920,    8*2048+ 987,   14*2048+1148,    0*2048+1355,
  41*2048+  13,    3*2048+ 261,   31*2048+ 422,    3*2048+ 572,   32*2048+ 709,   31*2048+ 792,   26*2048+ 853,   19*2048+ 882,    8*2048+ 883,    6*2048+ 938,   37*2048+1123,    3*2048+1190,    0*2048+1368,
   8*2048+ 392,   15*2048+ 451,    2*2048+ 548,   26*2048+ 601,    4*2048+ 608,   32*2048+ 668,   12*2048+ 728,   37*2048+ 793,    8*2048+ 901,   23*2048+ 980,   26*2048+1130,   32*2048+1290,    0*2048+1369,
  42*2048+  37,    4*2048+  91,   34*2048+ 134,    9*2048+ 183,   41*2048+ 560,    9*2048+ 573,   36*2048+ 745,    4*2048+ 782,   10*2048+ 829,    8*2048+1093,   28*2048+1184,   18*2048+1274,    0*2048+1370,
  21*2048+   1,   18*2048+   6,   32*2048+  38,   41*2048+ 477,   36*2048+ 590,   25*2048+ 626,   19*2048+ 673,   35*2048+ 751,   38*2048+ 758,   43*2048+ 854,   27*2048+ 861,   10*2048+1213,    0*2048+1371,
   2*2048+   2,   37*2048+  32,   30*2048+ 198,   20*2048+ 211,   45*2048+ 290,   41*2048+ 440,    1*2048+ 715,   22*2048+ 783,    4*2048+ 794,   27*2048+ 842,   20*2048+ 931,   41*2048+1291,    0*2048+1372,
  15*2048+  14,   19*2048+ 207,   12*2048+ 216,    4*2048+ 302,   24*2048+ 386,   45*2048+ 487,    9*2048+ 553,   43*2048+ 902,   10*2048+1052,    2*2048+1056,   22*2048+1082,    8*2048+1149,    0*2048+1373,
   4*2048+  56,   41*2048+ 175,    3*2048+ 423,   31*2048+ 584,    3*2048+ 734,   32*2048+ 871,   31*2048+ 955,   26*2048+1015,   19*2048+1045,    8*2048+1046,    6*2048+1101,   37*2048+1287,    0*2048+1386,
  33*2048+ 156,    8*2048+ 554,   15*2048+ 614,    2*2048+ 710,   26*2048+ 763,    4*2048+ 770,   32*2048+ 831,   12*2048+ 890,   37*2048+ 956,    8*2048+1063,   23*2048+1142,   26*2048+1292,    0*2048+1387,
  29*2048+  50,   19*2048+ 140,   42*2048+ 199,    4*2048+ 255,   34*2048+ 297,    9*2048+ 345,   41*2048+ 722,    9*2048+ 735,   36*2048+ 908,    4*2048+ 944,   10*2048+ 991,    8*2048+1256,    0*2048+1388,
  11*2048+  80,   21*2048+ 163,   18*2048+ 169,   32*2048+ 200,   41*2048+ 639,   36*2048+ 752,   25*2048+ 788,   19*2048+ 837,   35*2048+ 913,   38*2048+ 921,   43*2048+1016,   27*2048+1023,    0*2048+1389,
  42*2048+ 157,    2*2048+ 164,   37*2048+ 195,   30*2048+ 360,   20*2048+ 373,   45*2048+ 452,   41*2048+ 602,    1*2048+ 877,   22*2048+ 945,    4*2048+ 957,   27*2048+1004,   20*2048+1094,    0*2048+1390,
   9*2048+  15,   15*2048+ 176,   19*2048+ 369,   12*2048+ 379,    4*2048+ 464,   24*2048+ 549,   45*2048+ 651,    9*2048+ 716,   43*2048+1064,   10*2048+1214,    2*2048+1220,   22*2048+1244,    0*2048+1391,
  38*2048+ 153,    4*2048+ 218,   41*2048+ 337,    3*2048+ 585,   31*2048+ 746,    3*2048+ 896,   32*2048+1034,   31*2048+1117,   26*2048+1177,   19*2048+1208,    8*2048+1209,    6*2048+1263,    0*2048+1404,
  24*2048+   8,   27*2048+ 158,   33*2048+ 319,    8*2048+ 717,   15*2048+ 776,    2*2048+ 872,   26*2048+ 926,    4*2048+ 932,   32*2048+ 993,   12*2048+1053,   37*2048+1118,    8*2048+1226,    0*2048+1405,
   9*2048+ 122,   29*2048+ 213,   19*2048+ 303,   42*2048+ 361,    4*2048+ 417,   34*2048+ 459,    9*2048+ 507,   41*2048+ 884,    9*2048+ 897,   36*2048+1071,    4*2048+1106,   10*2048+1153,    0*2048+1406,
  11*2048+ 242,   21*2048+ 326,   18*2048+ 332,   32*2048+ 362,   41*2048+ 801,   36*2048+ 914,   25*2048+ 951,   19*2048+ 999,   35*2048+1076,   38*2048+1083,   43*2048+1178,   27*2048+1185,    0*2048+1407,
  42*2048+ 320,    2*2048+ 327,   37*2048+ 357,   30*2048+ 522,   20*2048+ 536,   45*2048+ 615,   41*2048+ 764,    1*2048+1040,   22*2048+1107,    4*2048+1119,   27*2048+1167,   20*2048+1257,    0*2048+1408,
  11*2048+  81,    3*2048+  86,   23*2048+ 111,    9*2048+ 177,   15*2048+ 338,   19*2048+ 531,   12*2048+ 542,    4*2048+ 627,   24*2048+ 711,   45*2048+ 813,    9*2048+ 878,   43*2048+1227,    0*2048+1409,
  27*2048+  43,   20*2048+  74,    9*2048+  75,    7*2048+ 129,   38*2048+ 315,    4*2048+ 381,   41*2048+ 500,    3*2048+ 747,   31*2048+ 909,    3*2048+1058,   32*2048+1197,   31*2048+1279,    0*2048+1422,
   9*2048+  92,   24*2048+ 171,   27*2048+ 321,   33*2048+ 482,    8*2048+ 879,   15*2048+ 939,    2*2048+1035,   26*2048+1089,    4*2048+1095,   32*2048+1155,   12*2048+1215,   37*2048+1280,    0*2048+1423,
  11*2048+  20,    9*2048+ 285,   29*2048+ 375,   19*2048+ 465,   42*2048+ 523,    4*2048+ 579,   34*2048+ 621,    9*2048+ 669,   41*2048+1047,    9*2048+1059,   36*2048+1233,    4*2048+1268,    0*2048+1424,
  44*2048+  44,   28*2048+  51,   11*2048+ 405,   21*2048+ 488,   18*2048+ 494,   32*2048+ 524,   41*2048+ 963,   36*2048+1077,   25*2048+1113,   19*2048+1161,   35*2048+1239,   38*2048+1245,    0*2048+1425,
  28*2048+  33,   21*2048+ 123,   42*2048+ 483,    2*2048+ 489,   37*2048+ 519,   30*2048+ 687,   20*2048+ 699,   45*2048+ 777,   41*2048+ 927,    1*2048+1203,   22*2048+1269,    4*2048+1281,    0*2048+1426,
  44*2048+  93,   11*2048+ 243,    3*2048+ 248,   23*2048+ 273,    9*2048+ 339,   15*2048+ 501,   19*2048+ 693,   12*2048+ 705,    4*2048+ 789,   24*2048+ 873,   45*2048+ 975,    9*2048+1041,    0*2048+1427,

   0*2048+   3,    0*2048+   9,    0*2048+1240,
   0*2048+  10,    0*2048+  16,    0*2048+1241,
   0*2048+  17,    0*2048+  22,    0*2048+1242,
   0*2048+  23,    0*2048+  26,    0*2048+1243,
   0*2048+  27,    0*2048+  31,    0*2048+1244,
   0*2048+  32,    0*2048+  35,    0*2048+1245,
   0*2048+  36,    0*2048+  40,    0*2048+1246,
   0*2048+  41,    0*2048+  46,    0*2048+1247,
   0*2048+  47,    0*2048+  51,    0*2048+1248,
   0*2048+  52,    0*2048+  56,    0*2048+1249,
   0*2048+  57,    0*2048+  62,    0*2048+1250,
   0*2048+  63,    0*2048+  68,    0*2048+1251,
   0*2048+  69,    0*2048+  74,    0*2048+1252,
   0*2048+  75,    0*2048+  80,    0*2048+1253,
   0*2048+  81,    0*2048+  85,    0*2048+1254,
   0*2048+  86,    0*2048+  89,    0*2048+1255,
   0*2048+  90,    0*2048+  95,    0*2048+1256,
   0*2048+  96,    0*2048+ 100,    0*2048+1257,
   0*2048+ 101,    0*2048+ 104,    0*2048+1258,
   0*2048+ 105,    0*2048+ 110,    0*2048+1259,
   0*2048+ 111,    0*2048+ 115,    0*2048+1260,
   0*2048+ 116,    0*2048+ 121,    0*2048+1261,
   0*2048+ 122,    0*2048+ 126,    0*2048+1262,
   0*2048+ 127,    0*2048+ 133,    0*2048+1263,
   0*2048+ 134,    0*2048+ 138,    0*2048+1264,
   0*2048+ 139,    0*2048+ 144,    0*2048+1265,
   0*2048+ 145,    0*2048+ 151,    0*2048+1266,
   0*2048+ 152,    0*2048+ 157,    0*2048+1267,
   0*2048+ 158,    0*2048+ 161,    0*2048+1268,
   0*2048+ 162,    0*2048+ 166,    0*2048+1269,
   0*2048+ 167,    0*2048+ 170,    0*2048+1270,
   0*2048+ 171,    0*2048+ 175,    0*2048+1271,
   0*2048+ 176,    0*2048+ 181,    0*2048+1272,
   0*2048+ 182,    0*2048+ 186,    0*2048+1273,
   0*2048+ 187,    0*2048+ 191,    0*2048+1274,
   0*2048+ 192,    0*2048+ 197,    0*2048+1275,
   0*2048+ 198,    0*2048+ 203,    0*2048+1276,
   0*2048+ 204,    0*2048+ 209,    0*2048+1277,
   0*2048+ 210,    0*2048+ 215,    0*2048+1278,
   0*2048+ 216,    0*2048+ 220,    0*2048+1279,
   0*2048+ 221,    0*2048+ 224,    0*2048+1280,
   0*2048+ 225,    0*2048+ 230,    0*2048+1281,
   0*2048+ 231,    0*2048+ 235,    0*2048+1282,
   0*2048+ 236,    0*2048+ 239,    0*2048+1283,
   0*2048+ 240,    0*2048+ 245,    0*2048+1284,
   0*2048+ 246,    0*2048+ 250,    0*2048+1285,
   0*2048+ 251,    0*2048+ 256,    0*2048+1286,
   0*2048+ 257,    0*2048+ 261,    0*2048+1287,
   0*2048+ 262,    0*2048+ 268,    0*2048+1288,
   0*2048+ 269,    0*2048+ 273,    0*2048+1289,
   0*2048+ 274,    0*2048+ 279,    0*2048+1290,
   0*2048+ 280,    0*2048+ 286,    0*2048+1291,
   0*2048+ 287,    0*2048+ 292,    0*2048+1292,
   0*2048+ 293,    0*2048+ 296,    0*2048+1293,
   0*2048+ 297,    0*2048+ 301,    0*2048+1294,
   0*2048+ 302,    0*2048+ 305,    0*2048+1295,
   0*2048+ 306,    0*2048+ 310,    0*2048+1296,
   0*2048+ 311,    0*2048+ 316,    0*2048+1297,
   0*2048+ 317,    0*2048+ 321,    0*2048+1298,
   0*2048+ 322,    0*2048+ 326,    0*2048+1299,
   0*2048+ 327,    0*2048+ 332,    0*2048+1300,
   0*2048+ 333,    0*2048+ 338,    0*2048+1301,
   0*2048+ 339,    0*2048+ 344,    0*2048+1302,
   0*2048+ 345,    0*2048+ 350,    0*2048+1303,
   0*2048+ 351,    0*2048+ 355,    0*2048+1304,
   0*2048+ 356,    0*2048+ 359,    0*2048+1305,
   0*2048+ 360,    0*2048+ 365,    0*2048+1306,
   0*2048+ 366,    0*2048+ 370,    0*2048+1307,
   0*2048+ 371,    0*2048+ 374,    0*2048+1308,
   0*2048+ 375,    0*2048+ 380,    0*2048+1309,
   0*2048+ 381,    0*2048+ 385,    0*2048+1310,
   0*2048+ 386,    0*2048+ 391,    0*2048+1311,
   0*2048+ 392,    0*2048+ 396,    0*2048+1312,
   0*2048+ 397,    0*2048+ 403,    0*2048+1313,
   0*2048+ 404,    0*2048+ 408,    0*2048+1314,
   0*2048+ 409,    0*2048+ 414,    0*2048+1315,
   0*2048+ 415,    0*2048+ 421,    0*2048+1316,
   0*2048+ 422,    0*2048+ 427,    0*2048+1317,
   0*2048+ 428,    0*2048+ 431,    0*2048+1318,
   0*2048+ 432,    0*2048+ 436,    0*2048+1319,
   0*2048+ 437,    0*2048+ 440,    0*2048+1320,
   0*2048+ 441,    0*2048+ 445,    0*2048+1321,
   0*2048+ 446,    0*2048+ 451,    0*2048+1322,
   0*2048+ 452,    0*2048+ 456,    0*2048+1323,
   0*2048+ 457,    0*2048+ 461,    0*2048+1324,
   0*2048+ 462,    0*2048+ 467,    0*2048+1325,
   0*2048+ 468,    0*2048+ 473,    0*2048+1326,
   0*2048+ 474,    0*2048+ 479,    0*2048+1327,
   0*2048+ 480,    0*2048+ 485,    0*2048+1328,
   0*2048+ 486,    0*2048+ 490,    0*2048+1329,
   0*2048+ 491,    0*2048+ 494,    0*2048+1330,
   0*2048+ 495,    0*2048+ 500,    0*2048+1331,
   0*2048+ 501,    0*2048+ 505,    0*2048+1332,
   0*2048+ 506,    0*2048+ 509,    0*2048+1333,
   0*2048+ 510,    0*2048+ 515,    0*2048+1334,
   0*2048+ 516,    0*2048+ 520,    0*2048+1335,
   0*2048+ 521,    0*2048+ 526,    0*2048+1336,
   0*2048+ 527,    0*2048+ 531,    0*2048+1337,
   0*2048+ 532,    0*2048+ 538,    0*2048+1338,
   0*2048+ 539,    0*2048+ 543,    0*2048+1339,
   0*2048+ 544,    0*2048+ 549,    0*2048+1340,
   0*2048+ 550,    0*2048+ 556,    0*2048+1341,
   0*2048+ 557,    0*2048+ 562,    0*2048+1342,
   0*2048+ 563,    0*2048+ 566,    0*2048+1343,
   0*2048+ 567,    0*2048+ 571,    0*2048+1344,
   0*2048+ 572,    0*2048+ 575,    0*2048+1345,
   0*2048+ 576,    0*2048+ 580,    0*2048+1346,
   0*2048+ 581,    0*2048+ 586,    0*2048+1347,
   0*2048+ 587,    0*2048+ 591,    0*2048+1348,
   0*2048+ 592,    0*2048+ 596,    0*2048+1349,
   0*2048+ 597,    0*2048+ 602,    0*2048+1350,
   0*2048+ 603,    0*2048+ 608,    0*2048+1351,
   0*2048+ 609,    0*2048+ 614,    0*2048+1352,
   0*2048+ 615,    0*2048+ 620,    0*2048+1353,
   0*2048+ 621,    0*2048+ 625,    0*2048+1354,
   0*2048+ 626,    0*2048+ 629,    0*2048+1355,
   0*2048+ 630,    0*2048+ 635,    0*2048+1356,
   0*2048+ 636,    0*2048+ 640,    0*2048+1357,
   0*2048+ 641,    0*2048+ 644,    0*2048+1358,
   0*2048+ 645,    0*2048+ 650,    0*2048+1359,
   0*2048+ 651,    0*2048+ 655,    0*2048+1360,
   0*2048+ 656,    0*2048+ 661,    0*2048+1361,
   0*2048+ 662,    0*2048+ 666,    0*2048+1362,
   0*2048+ 667,    0*2048+ 673,    0*2048+1363,
   0*2048+ 674,    0*2048+ 678,    0*2048+1364,
   0*2048+ 679,    0*2048+ 684,    0*2048+1365,
   0*2048+ 685,    0*2048+ 691,    0*2048+1366,
   0*2048+ 692,    0*2048+ 697,    0*2048+1367,
   0*2048+ 698,    0*2048+ 701,    0*2048+1368,
   0*2048+ 702,    0*2048+ 706,    0*2048+1369,
   0*2048+ 707,    0*2048+ 710,    0*2048+1370,
   0*2048+ 711,    0*2048+ 715,    0*2048+1371,
   0*2048+ 716,    0*2048+ 721,    0*2048+1372,
   0*2048+ 722,    0*2048+ 726,    0*2048+1373,
   0*2048+ 727,    0*2048+ 731,    0*2048+1374,
   0*2048+ 732,    0*2048+ 737,    0*2048+1375,
   0*2048+ 738,    0*2048+ 743,    0*2048+1376,
   0*2048+ 744,    0*2048+ 749,    0*2048+1377,
   0*2048+ 750,    0*2048+ 755,    0*2048+1378,
   0*2048+ 756,    0*2048+ 760,    0*2048+1379,
   0*2048+ 761,    0*2048+ 764,    0*2048+1380,
   0*2048+ 765,    0*2048+ 770,    0*2048+1381,
   0*2048+ 771,    0*2048+ 775,    0*2048+1382,
   0*2048+ 776,    0*2048+ 779,    0*2048+1383,
   0*2048+ 780,    0*2048+ 785,    0*2048+1384,
   0*2048+ 786,    0*2048+ 790,    0*2048+1385,
   0*2048+ 791,    0*2048+ 796,    0*2048+1386,
   0*2048+ 797,    0*2048+ 801,    0*2048+1387,
   0*2048+ 802,    0*2048+ 808,    0*2048+1388,
   0*2048+ 809,    0*2048+ 813,    0*2048+1389,
   0*2048+ 814,    0*2048+ 819,    0*2048+1390,
   0*2048+ 820,    0*2048+ 826,    0*2048+1391,
   0*2048+ 827,    0*2048+ 832,    0*2048+1392,
   0*2048+ 833,    0*2048+ 836,    0*2048+1393,
   0*2048+ 837,    0*2048+ 841,    0*2048+1394,
   0*2048+ 842,    0*2048+ 845,    0*2048+1395,
   0*2048+ 846,    0*2048+ 850,    0*2048+1396,
   0*2048+ 851,    0*2048+ 856,    0*2048+1397,
   0*2048+ 857,    0*2048+ 861,    0*2048+1398,
   0*2048+ 862,    0*2048+ 866,    0*2048+1399,
   0*2048+ 867,    0*2048+ 872,    0*2048+1400,
   0*2048+ 873,    0*2048+ 878,    0*2048+1401,
   0*2048+ 879,    0*2048+ 884,    0*2048+1402,
   0*2048+ 885,    0*2048+ 890,    0*2048+1403,
   0*2048+ 891,    0*2048+ 895,    0*2048+1404,
   0*2048+ 896,    0*2048+ 899,    0*2048+1405,
   0*2048+ 900,    0*2048+ 905,    0*2048+1406,
   0*2048+ 906,    0*2048+ 910,    0*2048+1407,
   0*2048+ 911,    0*2048+ 914,    0*2048+1408,
   0*2048+ 915,    0*2048+ 920,    0*2048+1409,
   0*2048+ 921,    0*2048+ 925,    0*2048+1410,
   0*2048+ 926,    0*2048+ 931,    0*2048+1411,
   0*2048+ 932,    0*2048+ 936,    0*2048+1412,
   0*2048+ 937,    0*2048+ 943,    0*2048+1413,
   0*2048+ 944,    0*2048+ 948,    0*2048+1414,
   0*2048+ 949,    0*2048+ 954,    0*2048+1415,
   0*2048+ 955,    0*2048+ 961,    0*2048+1416,
   0*2048+ 962,    0*2048+ 967,    0*2048+1417,
   0*2048+ 968,    0*2048+ 971,    0*2048+1418,
   0*2048+ 972,    0*2048+ 976,    0*2048+1419,
   0*2048+ 977,    0*2048+ 980,    0*2048+1420,
   0*2048+ 981,    0*2048+ 985,    0*2048+1421,
   0*2048+ 986,    0*2048+ 991,    0*2048+1422,
   0*2048+ 992,    0*2048+ 996,    0*2048+1423,
   0*2048+ 997,    0*2048+1001,    0*2048+1424,
   0*2048+1002,    0*2048+1007,    0*2048+1425,
   0*2048+1008,    0*2048+1013,    0*2048+1426,
   0*2048+1014,    0*2048+1019,    0*2048+1427,
   0*2048+1020,    0*2048+1025,    0*2048+1428,
   0*2048+1026,    0*2048+1030,    0*2048+1429,
   0*2048+1031,    0*2048+1034,    0*2048+1430,
   0*2048+1035,    0*2048+1040,    0*2048+1431,
   0*2048+1041,    0*2048+1045,    0*2048+1432,
   0*2048+1046,    0*2048+1049,    0*2048+1433,
   0*2048+1050,    0*2048+1055,    0*2048+1434,
   0*2048+1056,    0*2048+1060,    0*2048+1435,
   0*2048+1061,    0*2048+1066,    0*2048+1436,
   0*2048+1067,    0*2048+1071,    0*2048+1437,
   0*2048+1072,    0*2048+1078,    0*2048+1438,
   1*2048+   4,    0*2048+1079,    0*2048+1439,
   0*2048+   0,   20*2048+ 247,   34*2048+ 723,    0*2048+1085,
   0*2048+   5,   14*2048+ 298,    0*2048+ 357,    0*2048+1086,
   0*2048+  13,    1*2048+  64,   33*2048+ 507,    0*2048+1087,
   0*2048+  19,   17*2048+ 211,    5*2048+ 853,    0*2048+1088,
   0*2048+  24,   22*2048+ 119,   19*2048+ 270,    0*2048+1089,
   0*2048+  28,    1*2048+ 487,   29*2048+ 669,    0*2048+1090,
   0*2048+  33,   20*2048+ 264,    7*2048+ 362,    0*2048+1091,
   0*2048+  37,   39*2048+ 107,   11*2048+ 226,    0*2048+1092,
  23*2048+  34,    0*2048+  42,   15*2048+ 433,    0*2048+1093,
   0*2048+  48,   23*2048+ 177,   39*2048+ 416,    0*2048+1094,
   0*2048+  53,   34*2048+ 367,   19*2048+ 453,    0*2048+1095,
   0*2048+  58,   44*2048+ 728,   24*2048+1057,    0*2048+1096,
   0*2048+  65,   15*2048+ 153,    3*2048+ 886,    0*2048+1097,
   0*2048+  70,    5*2048+ 307,   29*2048+1015,    0*2048+1098,
  37*2048+  59,    0*2048+  76,   17*2048+ 271,    0*2048+1099,
   0*2048+ 135,   20*2048+ 382,   34*2048+ 858,    0*2048+1105,
   0*2048+ 140,   14*2048+ 434,    0*2048+ 493,    0*2048+1106,
   0*2048+ 148,    1*2048+ 199,   33*2048+ 642,    0*2048+1107,
   0*2048+ 155,   17*2048+ 346,    5*2048+ 988,    0*2048+1108,
   0*2048+ 159,   22*2048+ 254,   19*2048+ 405,    0*2048+1109,
   0*2048+ 163,    1*2048+ 622,   29*2048+ 804,    0*2048+1110,
   0*2048+ 168,   20*2048+ 399,    7*2048+ 497,    0*2048+1111,
   0*2048+ 172,   39*2048+ 243,   11*2048+ 363,    0*2048+1112,
  23*2048+ 169,    0*2048+ 178,   15*2048+ 568,    0*2048+1113,
   0*2048+ 183,   23*2048+ 312,   39*2048+ 551,    0*2048+1114,
   0*2048+ 188,   34*2048+ 503,   19*2048+ 588,    0*2048+1115,
  25*2048+ 113,    0*2048+ 193,   44*2048+ 863,    0*2048+1116,
   0*2048+ 200,   15*2048+ 288,    3*2048+1021,    0*2048+1117,
  30*2048+  71,    0*2048+ 206,    5*2048+ 442,    0*2048+1118,
  37*2048+ 194,    0*2048+ 212,   17*2048+ 406,    0*2048+1119,
   0*2048+ 272,   20*2048+ 517,   34*2048+ 993,    0*2048+1125,
   0*2048+ 275,   14*2048+ 569,    0*2048+ 628,    0*2048+1126,
   0*2048+ 283,    1*2048+ 335,   33*2048+ 777,    0*2048+1127,
   6*2048+  44,    0*2048+ 290,   17*2048+ 482,    0*2048+1128,
   0*2048+ 294,   22*2048+ 389,   19*2048+ 540,    0*2048+1129,
   0*2048+ 299,    1*2048+ 758,   29*2048+ 939,    0*2048+1130,
   0*2048+ 303,   20*2048+ 534,    7*2048+ 632,    0*2048+1131,
   0*2048+ 308,   39*2048+ 378,   11*2048+ 498,    0*2048+1132,
  23*2048+ 304,    0*2048+ 313,   15*2048+ 703,    0*2048+1133,
   0*2048+ 318,   23*2048+ 447,   39*2048+ 686,    0*2048+1134,
   0*2048+ 323,   34*2048+ 638,   19*2048+ 724,    0*2048+1135,
  25*2048+ 249,    0*2048+ 329,   44*2048+ 999,    0*2048+1136,
   4*2048+  77,    0*2048+ 336,   15*2048+ 423,    0*2048+1137,
  30*2048+ 207,    0*2048+ 342,    5*2048+ 578,    0*2048+1138,
  37*2048+ 330,    0*2048+ 347,   17*2048+ 541,    0*2048+1139,
  35*2048+  49,    0*2048+ 407,   20*2048+ 652,    0*2048+1145,
   0*2048+ 411,   14*2048+ 704,    0*2048+ 763,    0*2048+1146,
   0*2048+ 419,    1*2048+ 470,   33*2048+ 912,    0*2048+1147,
   6*2048+ 180,    0*2048+ 425,   17*2048+ 617,    0*2048+1148,
   0*2048+ 429,   22*2048+ 525,   19*2048+ 675,    0*2048+1149,
   0*2048+ 435,    1*2048+ 893,   29*2048+1074,    0*2048+1150,
   0*2048+ 438,   20*2048+ 671,    7*2048+ 768,    0*2048+1151,
   0*2048+ 443,   39*2048+ 513,   11*2048+ 633,    0*2048+1152,
  23*2048+ 439,    0*2048+ 448,   15*2048+ 838,    0*2048+1153,
   0*2048+ 454,   23*2048+ 582,   39*2048+ 821,    0*2048+1154,
   0*2048+ 458,   34*2048+ 774,   19*2048+ 859,    0*2048+1155,
  45*2048+  55,   25*2048+ 384,    0*2048+ 464,    0*2048+1156,
   4*2048+ 213,    0*2048+ 471,   15*2048+ 558,    0*2048+1157,
  30*2048+ 343,    0*2048+ 477,    5*2048+ 713,    0*2048+1158,
  37*2048+ 465,    0*2048+ 483,   17*2048+ 676,    0*2048+1159,
  35*2048+ 184,    0*2048+ 542,   20*2048+ 787,    0*2048+1165,
   0*2048+ 547,   14*2048+ 839,    0*2048+ 898,    0*2048+1166,
   0*2048+ 554,    1*2048+ 606,   33*2048+1047,    0*2048+1167,
   6*2048+ 315,    0*2048+ 560,   17*2048+ 752,    0*2048+1168,
   0*2048+ 564,   22*2048+ 660,   19*2048+ 810,    0*2048+1169,
  30*2048+ 130,    0*2048+ 570,    1*2048+1029,    0*2048+1170,
   0*2048+ 573,   20*2048+ 806,    7*2048+ 903,    0*2048+1171,
   0*2048+ 579,   39*2048+ 649,   11*2048+ 769,    0*2048+1172,
  23*2048+ 574,    0*2048+ 583,   15*2048+ 973,    0*2048+1173,
   0*2048+ 589,   23*2048+ 717,   39*2048+ 957,    0*2048+1174,
   0*2048+ 593,   34*2048+ 909,   19*2048+ 994,    0*2048+1175,
  45*2048+ 190,   25*2048+ 519,    0*2048+ 599,    0*2048+1176,
   4*2048+ 348,    0*2048+ 607,   15*2048+ 694,    0*2048+1177,
  30*2048+ 478,    0*2048+ 612,    5*2048+ 848,    0*2048+1178,
  37*2048+ 600,    0*2048+ 618,   17*2048+ 811,    0*2048+1179,
  35*2048+ 319,    0*2048+ 677,   20*2048+ 922,    0*2048+1185,
   0*2048+ 683,   14*2048+ 974,    0*2048+1033,    0*2048+1186,
  34*2048+ 102,    0*2048+ 689,    1*2048+ 741,    0*2048+1187,
   6*2048+ 450,    0*2048+ 696,   17*2048+ 888,    0*2048+1188,
   0*2048+ 699,   22*2048+ 795,   19*2048+ 945,    0*2048+1189,
   2*2048+  84,   30*2048+ 267,    0*2048+ 705,    0*2048+1190,
   0*2048+ 708,   20*2048+ 941,    7*2048+1038,    0*2048+1191,
   0*2048+ 714,   39*2048+ 784,   11*2048+ 904,    0*2048+1192,
  16*2048+  29,   23*2048+ 709,    0*2048+ 718,    0*2048+1193,
  40*2048+  15,    0*2048+ 725,   23*2048+ 854,    0*2048+1194,
  20*2048+  50,    0*2048+ 729,   34*2048+1044,    0*2048+1195,
  45*2048+ 325,   25*2048+ 654,    0*2048+ 734,    0*2048+1196,
   4*2048+ 484,    0*2048+ 742,   15*2048+ 829,    0*2048+1197,
  30*2048+ 613,    0*2048+ 747,    5*2048+ 983,    0*2048+1198,
  37*2048+ 735,    0*2048+ 753,   17*2048+ 946,    0*2048+1199,
  35*2048+ 455,    0*2048+ 812,   20*2048+1058,    0*2048+1205,
  15*2048+  30,    1*2048+  88,    0*2048+ 818,    0*2048+1206,
  34*2048+ 237,    0*2048+ 824,    1*2048+ 876,    0*2048+1207,
   6*2048+ 585,    0*2048+ 831,   17*2048+1023,    0*2048+1208,
  20*2048+   1,    0*2048+ 835,   22*2048+ 930,    0*2048+1209,
   2*2048+ 219,   30*2048+ 402,    0*2048+ 840,    0*2048+1210,
   8*2048+  93,    0*2048+ 843,   20*2048+1076,    0*2048+1211,
   0*2048+ 849,   39*2048+ 919,   11*2048+1039,    0*2048+1212,
  16*2048+ 164,   23*2048+ 844,    0*2048+ 855,    0*2048+1213,
  40*2048+ 150,    0*2048+ 860,   23*2048+ 989,    0*2048+1214,
  35*2048+  99,   20*2048+ 185,    0*2048+ 864,    0*2048+1215,
  45*2048+ 460,   25*2048+ 789,    0*2048+ 869,    0*2048+1216,
   4*2048+ 619,    0*2048+ 877,   15*2048+ 964,    0*2048+1217,
   6*2048+  39,   30*2048+ 748,    0*2048+ 882,    0*2048+1218,
  18*2048+   2,   37*2048+ 870,    0*2048+ 889,    0*2048+1219,
  21*2048+ 114,   35*2048+ 590,    0*2048+ 947,    0*2048+1225,
  15*2048+ 165,    1*2048+ 223,    0*2048+ 953,    0*2048+1226,
  34*2048+ 373,    0*2048+ 960,    1*2048+1011,    0*2048+1227,
  18*2048+  79,    6*2048+ 720,    0*2048+ 966,    0*2048+1228,
  20*2048+ 136,    0*2048+ 970,   22*2048+1065,    0*2048+1229,
   2*2048+ 354,   30*2048+ 537,    0*2048+ 975,    0*2048+1230,
  21*2048+ 132,    8*2048+ 229,    0*2048+ 978,    0*2048+1231,
  12*2048+  94,    0*2048+ 984,   39*2048+1054,    0*2048+1232,
  16*2048+ 300,   23*2048+ 979,    0*2048+ 990,    0*2048+1233,
  24*2048+  45,   40*2048+ 285,    0*2048+ 995,    0*2048+1234,
  35*2048+ 234,   20*2048+ 320,    0*2048+1000,    0*2048+1235,
  45*2048+ 595,   25*2048+ 924,    0*2048+1005,    0*2048+1236,
  16*2048+  21,    4*2048+ 754,    0*2048+1012,    0*2048+1237,
   6*2048+ 174,   30*2048+ 883,    0*2048+1018,    0*2048+1238,
  18*2048+ 137,   37*2048+1006,    0*2048+1024,    0*2048+1239,
   0*2048+ 106,   25*2048+ 241,   20*2048+ 328,    5*2048+ 334,    3*2048+ 604,   31*2048+ 834,   25*2048+ 852,   11*2048+1003,    0*2048+1080,
   0*2048+ 112,   24*2048+ 117,   29*2048+ 410,   15*2048+ 481,   31*2048+ 693,   12*2048+ 772,   28*2048+ 798,   11*2048+ 799,    0*2048+1081,
   0*2048+ 118,   12*2048+ 205,    1*2048+ 372,   18*2048+ 502,   28*2048+ 545,   17*2048+ 577,    4*2048+ 680,   15*2048+1027,    0*2048+1082,
  14*2048+  11,    0*2048+ 123,   22*2048+ 263,   23*2048+ 361,    5*2048+ 492,   22*2048+ 646,   26*2048+ 668,   17*2048+ 956,    0*2048+1083,
  31*2048+  12,   10*2048+  18,    0*2048+ 128,    6*2048+ 340,   32*2048+ 522,   25*2048+ 757,   23*2048+ 766,    5*2048+ 998,    0*2048+1084,
  12*2048+  60,    0*2048+ 242,   25*2048+ 376,   20*2048+ 463,    5*2048+ 469,    3*2048+ 739,   31*2048+ 969,   25*2048+ 987,    0*2048+1100,
   0*2048+ 248,   24*2048+ 252,   29*2048+ 546,   15*2048+ 616,   31*2048+ 828,   12*2048+ 907,   28*2048+ 933,   11*2048+ 934,    0*2048+1101,
  16*2048+  82,    0*2048+ 253,   12*2048+ 341,    1*2048+ 508,   18*2048+ 637,   28*2048+ 681,   17*2048+ 712,    4*2048+ 815,    0*2048+1102,
  18*2048+  14,   14*2048+ 146,    0*2048+ 258,   22*2048+ 398,   23*2048+ 496,    5*2048+ 627,   22*2048+ 781,   26*2048+ 803,    0*2048+1103,
   6*2048+  54,   31*2048+ 147,   10*2048+ 154,    0*2048+ 265,    6*2048+ 475,   32*2048+ 657,   25*2048+ 892,   23*2048+ 901,    0*2048+1104,
  32*2048+  25,   26*2048+  43,   12*2048+ 195,    0*2048+ 377,   25*2048+ 511,   20*2048+ 598,    5*2048+ 605,    3*2048+ 874,    0*2048+1120,
   0*2048+ 383,   24*2048+ 387,   29*2048+ 682,   15*2048+ 751,   31*2048+ 963,   12*2048+1042,   28*2048+1068,   11*2048+1069,    0*2048+1121,
  16*2048+ 217,    0*2048+ 388,   12*2048+ 476,    1*2048+ 643,   18*2048+ 773,   28*2048+ 816,   17*2048+ 847,    4*2048+ 950,    0*2048+1122,
  18*2048+ 149,   14*2048+ 281,    0*2048+ 393,   22*2048+ 533,   23*2048+ 631,    5*2048+ 762,   22*2048+ 916,   26*2048+ 938,    0*2048+1123,
   6*2048+ 189,   31*2048+ 282,   10*2048+ 289,    0*2048+ 400,    6*2048+ 610,   32*2048+ 792,   25*2048+1028,   23*2048+1036,    0*2048+1124,
  32*2048+ 160,   26*2048+ 179,   12*2048+ 331,    0*2048+ 512,   25*2048+ 647,   20*2048+ 733,    5*2048+ 740,    3*2048+1009,    0*2048+1140,
  32*2048+  20,   13*2048+  97,   29*2048+ 124,   12*2048+ 125,    0*2048+ 518,   24*2048+ 523,   29*2048+ 817,   15*2048+ 887,    0*2048+1141,
   5*2048+   6,   16*2048+ 352,    0*2048+ 524,   12*2048+ 611,    1*2048+ 778,   18*2048+ 908,   28*2048+ 951,   17*2048+ 982,    0*2048+1142,
  18*2048+ 284,   14*2048+ 417,    0*2048+ 528,   22*2048+ 670,   23*2048+ 767,    5*2048+ 897,   22*2048+1051,   26*2048+1073,    0*2048+1143,
  26*2048+  83,   24*2048+  91,    6*2048+ 324,   31*2048+ 418,   10*2048+ 424,    0*2048+ 535,    6*2048+ 745,   32*2048+ 927,    0*2048+1144,
   4*2048+  66,   32*2048+ 295,   26*2048+ 314,   12*2048+ 466,    0*2048+ 648,   25*2048+ 782,   20*2048+ 868,    5*2048+ 875,    0*2048+1160,
  32*2048+ 156,   13*2048+ 232,   29*2048+ 259,   12*2048+ 260,    0*2048+ 653,   24*2048+ 658,   29*2048+ 952,   15*2048+1022,    0*2048+1161,
  29*2048+   7,   18*2048+  38,    5*2048+ 141,   16*2048+ 488,    0*2048+ 659,   12*2048+ 746,    1*2048+ 913,   18*2048+1043,    0*2048+1162,
  23*2048+ 108,   27*2048+ 129,   18*2048+ 420,   14*2048+ 552,    0*2048+ 663,   22*2048+ 805,   23*2048+ 902,    5*2048+1032,    0*2048+1163,
  26*2048+ 218,   24*2048+ 227,    6*2048+ 459,   31*2048+ 553,   10*2048+ 559,    0*2048+ 672,    6*2048+ 880,   32*2048+1062,    0*2048+1164,
   4*2048+ 201,   32*2048+ 430,   26*2048+ 449,   12*2048+ 601,    0*2048+ 783,   25*2048+ 917,   20*2048+1004,    5*2048+1010,    0*2048+1180,
  30*2048+   8,   16*2048+  78,   32*2048+ 291,   13*2048+ 368,   29*2048+ 394,   12*2048+ 395,    0*2048+ 788,   24*2048+ 793,    0*2048+1181,
  19*2048+  98,   29*2048+ 142,   18*2048+ 173,    5*2048+ 276,   16*2048+ 623,    0*2048+ 794,   12*2048+ 881,    1*2048+1048,    0*2048+1182,
   6*2048+  87,   23*2048+ 244,   27*2048+ 266,   18*2048+ 555,   14*2048+ 687,    0*2048+ 800,   22*2048+ 940,   23*2048+1037,    0*2048+1183,
  33*2048+ 120,   26*2048+ 353,   24*2048+ 364,    6*2048+ 594,   31*2048+ 688,   10*2048+ 695,    0*2048+ 807,    6*2048+1016,    0*2048+1184,
  21*2048+  61,    6*2048+  67,    4*2048+ 337,   32*2048+ 565,   26*2048+ 584,   12*2048+ 736,    0*2048+ 918,   25*2048+1052,    0*2048+1200,
  30*2048+ 143,   16*2048+ 214,   32*2048+ 426,   13*2048+ 504,   29*2048+ 529,   12*2048+ 530,    0*2048+ 923,   24*2048+ 928,    0*2048+1201,
   2*2048+ 103,   19*2048+ 233,   29*2048+ 277,   18*2048+ 309,    5*2048+ 412,   16*2048+ 759,    0*2048+ 929,   12*2048+1017,    0*2048+1202,
  24*2048+  92,    6*2048+ 222,   23*2048+ 379,   27*2048+ 401,   18*2048+ 690,   14*2048+ 822,    0*2048+ 935,   22*2048+1075,    0*2048+1203,
   7*2048+  72,   33*2048+ 255,   26*2048+ 489,   24*2048+ 499,    6*2048+ 730,   31*2048+ 823,   10*2048+ 830,    0*2048+ 942,    0*2048+1204,
  26*2048+ 109,   21*2048+ 196,    6*2048+ 202,    4*2048+ 472,   32*2048+ 700,   26*2048+ 719,   12*2048+ 871,    0*2048+1053,    0*2048+1220,
  30*2048+ 278,   16*2048+ 349,   32*2048+ 561,   13*2048+ 639,   29*2048+ 664,   12*2048+ 665,    0*2048+1059,   24*2048+1063,    0*2048+1221,
  13*2048+  73,    2*2048+ 238,   19*2048+ 369,   29*2048+ 413,   18*2048+ 444,    5*2048+ 548,   16*2048+ 894,    0*2048+1064,    0*2048+1222,
  23*2048+ 131,   24*2048+ 228,    6*2048+ 358,   23*2048+ 514,   27*2048+ 536,   18*2048+ 825,   14*2048+ 958,    0*2048+1070,    0*2048+1223,
   7*2048+ 208,   33*2048+ 390,   26*2048+ 624,   24*2048+ 634,    6*2048+ 865,   31*2048+ 959,   10*2048+ 965,    0*2048+1077,    0*2048+1224,

   0*2048+   9,    0*2048+  20,    0*2048+1800,
   0*2048+  21,    0*2048+  31,    0*2048+1801,
   0*2048+  32,    0*2048+  42,    0*2048+1802,
   0*2048+  43,    0*2048+  53,    0*2048+1803,
   0*2048+  54,    0*2048+  64,    0*2048+1804,
   0*2048+  65,    0*2048+  75,    0*2048+1805,
   0*2048+  76,    0*2048+  86,    0*2048+1806,
   0*2048+  87,    0*2048+  97,    0*2048+1807,
   0*2048+  98,    0*2048+ 108,    0*2048+1808,
   0*2048+ 109,    0*2048+ 119,    0*2048+1809,
   0*2048+ 120,    0*2048+ 130,    0*2048+1810,
   0*2048+ 131,    0*2048+ 141,    0*2048+1811,
   0*2048+ 142,    0*2048+ 152,    0*2048+1812,
   0*2048+ 153,    0*2048+ 163,    0*2048+1813,
   0*2048+ 164,    0*2048+ 174,    0*2048+1814,
   0*2048+ 175,    0*2048+ 185,    0*2048+1815,
   0*2048+ 186,    0*2048+ 196,    0*2048+1816,
   0*2048+ 197,    0*2048+ 207,    0*2048+1817,
   0*2048+ 208,    0*2048+ 218,    0*2048+1818,
   0*2048+ 219,    0*2048+ 229,    0*2048+1819,
   0*2048+ 230,    0*2048+ 240,    0*2048+1820,
   0*2048+ 241,    0*2048+ 251,    0*2048+1821,
   0*2048+ 252,    0*2048+ 262,    0*2048+1822,
   0*2048+ 263,    0*2048+ 273,    0*2048+1823,
   0*2048+ 274,    0*2048+ 284,    0*2048+1824,
   0*2048+ 285,    0*2048+ 295,    0*2048+1825,
   0*2048+ 296,    0*2048+ 306,    0*2048+1826,
   0*2048+ 307,    0*2048+ 317,    0*2048+1827,
   0*2048+ 318,    0*2048+ 328,    0*2048+1828,
   0*2048+ 329,    0*2048+ 339,    0*2048+1829,
   0*2048+ 340,    0*2048+ 350,    0*2048+1830,
   0*2048+ 351,    0*2048+ 361,    0*2048+1831,
   0*2048+ 362,    0*2048+ 372,    0*2048+1832,
   0*2048+ 373,    0*2048+ 383,    0*2048+1833,
   0*2048+ 384,    0*2048+ 394,    0*2048+1834,
   0*2048+ 395,    0*2048+ 405,    0*2048+1835,
   0*2048+ 406,    0*2048+ 416,    0*2048+1836,
   0*2048+ 417,    0*2048+ 427,    0*2048+1837,
   0*2048+ 428,    0*2048+ 438,    0*2048+1838,
   0*2048+ 439,    0*2048+ 449,    0*2048+1839,
   0*2048+ 450,    0*2048+ 460,    0*2048+1840,
   0*2048+ 461,    0*2048+ 471,    0*2048+1841,
   0*2048+ 472,    0*2048+ 482,    0*2048+1842,
   0*2048+ 483,    0*2048+ 493,    0*2048+1843,
   0*2048+ 494,    0*2048+ 504,    0*2048+1844,
   0*2048+ 505,    0*2048+ 515,    0*2048+1845,
   0*2048+ 516,    0*2048+ 526,    0*2048+1846,
   0*2048+ 527,    0*2048+ 537,    0*2048+1847,
   0*2048+ 538,    0*2048+ 548,    0*2048+1848,
   0*2048+ 549,    0*2048+ 559,    0*2048+1849,
   0*2048+ 560,    0*2048+ 570,    0*2048+1850,
   0*2048+ 571,    0*2048+ 581,    0*2048+1851,
   0*2048+ 582,    0*2048+ 592,    0*2048+1852,
   0*2048+ 593,    0*2048+ 603,    0*2048+1853,
   0*2048+ 604,    0*2048+ 614,    0*2048+1854,
   0*2048+ 615,    0*2048+ 625,    0*2048+1855,
   0*2048+ 626,    0*2048+ 636,    0*2048+1856,
   0*2048+ 637,    0*2048+ 647,    0*2048+1857,
   0*2048+ 648,    0*2048+ 658,    0*2048+1858,
   0*2048+ 659,    0*2048+ 669,    0*2048+1859,
   0*2048+ 670,    0*2048+ 680,    0*2048+1860,
   0*2048+ 681,    0*2048+ 691,    0*2048+1861,
   0*2048+ 692,    0*2048+ 702,    0*2048+1862,
   0*2048+ 703,    0*2048+ 713,    0*2048+1863,
   0*2048+ 714,    0*2048+ 724,    0*2048+1864,
   0*2048+ 725,    0*2048+ 735,    0*2048+1865,
   0*2048+ 736,    0*2048+ 746,    0*2048+1866,
   0*2048+ 747,    0*2048+ 757,    0*2048+1867,
   0*2048+ 758,    0*2048+ 768,    0*2048+1868,
   0*2048+ 769,    0*2048+ 779,    0*2048+1869,
   0*2048+ 780,    0*2048+ 790,    0*2048+1870,
   0*2048+ 791,    0*2048+ 801,    0*2048+1871,
   0*2048+ 802,    0*2048+ 812,    0*2048+1872,
   0*2048+ 813,    0*2048+ 823,    0*2048+1873,
   0*2048+ 824,    0*2048+ 834,    0*2048+1874,
   0*2048+ 835,    0*2048+ 845,    0*2048+1875,
   0*2048+ 846,    0*2048+ 856,    0*2048+1876,
   0*2048+ 857,    0*2048+ 867,    0*2048+1877,
   0*2048+ 868,    0*2048+ 878,    0*2048+1878,
   0*2048+ 879,    0*2048+ 889,    0*2048+1879,
   0*2048+ 890,    0*2048+ 900,    0*2048+1880,
   0*2048+ 901,    0*2048+ 911,    0*2048+1881,
   0*2048+ 912,    0*2048+ 922,    0*2048+1882,
   0*2048+ 923,    0*2048+ 933,    0*2048+1883,
   0*2048+ 934,    0*2048+ 944,    0*2048+1884,
   0*2048+ 945,    0*2048+ 955,    0*2048+1885,
   0*2048+ 956,    0*2048+ 966,    0*2048+1886,
   0*2048+ 967,    0*2048+ 977,    0*2048+1887,
   0*2048+ 978,    0*2048+ 988,    0*2048+1888,
   0*2048+ 989,    0*2048+ 999,    0*2048+1889,
   0*2048+1000,    0*2048+1010,    0*2048+1890,
   0*2048+1011,    0*2048+1021,    0*2048+1891,
   0*2048+1022,    0*2048+1032,    0*2048+1892,
   0*2048+1033,    0*2048+1043,    0*2048+1893,
   0*2048+1044,    0*2048+1054,    0*2048+1894,
   0*2048+1055,    0*2048+1065,    0*2048+1895,
   0*2048+1066,    0*2048+1076,    0*2048+1896,
   0*2048+1077,    0*2048+1087,    0*2048+1897,
   0*2048+1088,    0*2048+1098,    0*2048+1898,
   0*2048+1099,    0*2048+1109,    0*2048+1899,
   0*2048+1110,    0*2048+1120,    0*2048+1900,
   0*2048+1121,    0*2048+1131,    0*2048+1901,
   0*2048+1132,    0*2048+1142,    0*2048+1902,
   0*2048+1143,    0*2048+1153,    0*2048+1903,
   0*2048+1154,    0*2048+1164,    0*2048+1904,
   0*2048+1165,    0*2048+1175,    0*2048+1905,
   0*2048+1176,    0*2048+1186,    0*2048+1906,
   0*2048+1187,    0*2048+1197,    0*2048+1907,
   0*2048+1198,    0*2048+1208,    0*2048+1908,
   0*2048+1209,    0*2048+1219,    0*2048+1909,
   0*2048+1220,    0*2048+1230,    0*2048+1910,
   0*2048+1231,    0*2048+1241,    0*2048+1911,
   0*2048+1242,    0*2048+1252,    0*2048+1912,
   0*2048+1253,    0*2048+1263,    0*2048+1913,
   0*2048+1264,    0*2048+1274,    0*2048+1914,
   0*2048+1275,    0*2048+1285,    0*2048+1915,
   0*2048+1286,    0*2048+1296,    0*2048+1916,
   0*2048+1297,    0*2048+1307,    0*2048+1917,
   0*2048+1308,    0*2048+1318,    0*2048+1918,
   0*2048+1319,    0*2048+1329,    0*2048+1919,
   0*2048+1330,    0*2048+1340,    0*2048+1920,
   0*2048+1341,    0*2048+1351,    0*2048+1921,
   0*2048+1352,    0*2048+1362,    0*2048+1922,
   0*2048+1363,    0*2048+1373,    0*2048+1923,
   0*2048+1374,    0*2048+1384,    0*2048+1924,
   0*2048+1385,    0*2048+1395,    0*2048+1925,
   0*2048+1396,    0*2048+1406,    0*2048+1926,
   0*2048+1407,    0*2048+1417,    0*2048+1927,
   0*2048+1418,    0*2048+1428,    0*2048+1928,
   0*2048+1429,    0*2048+1439,    0*2048+1929,
   0*2048+1440,    0*2048+1450,    0*2048+1930,
   0*2048+1451,    0*2048+1461,    0*2048+1931,
   0*2048+1462,    0*2048+1472,    0*2048+1932,
   0*2048+1473,    0*2048+1483,    0*2048+1933,
   0*2048+1484,    0*2048+1494,    0*2048+1934,
   0*2048+1495,    0*2048+1505,    0*2048+1935,
   0*2048+1506,    0*2048+1516,    0*2048+1936,
   0*2048+1517,    0*2048+1527,    0*2048+1937,
   0*2048+1528,    0*2048+1538,    0*2048+1938,
   0*2048+1539,    0*2048+1549,    0*2048+1939,
   0*2048+1550,    0*2048+1560,    0*2048+1940,
   0*2048+1561,    0*2048+1571,    0*2048+1941,
   0*2048+1572,    0*2048+1582,    0*2048+1942,
   1*2048+  10,    0*2048+1583,    0*2048+1943,
   0*2048+   0,   15*2048+  11,   18*2048+ 671,    0*2048+1593,
   0*2048+  12,   10*2048+ 231,    9*2048+ 924,    0*2048+1594,
   0*2048+  22,   17*2048+ 594,   25*2048+1177,    0*2048+1595,
   0*2048+  35,    7*2048+ 540,   27*2048+ 913,    0*2048+1596,
   0*2048+  44,   42*2048+ 154,   41*2048+ 892,    0*2048+1597,
   0*2048+  56,   12*2048+  57,   41*2048+1366,    0*2048+1598,
   0*2048+  66,   26*2048+ 463,   13*2048+ 704,    0*2048+1599,
   0*2048+  78,    6*2048+1012,   29*2048+1276,    0*2048+1600,
   0*2048+  88,   39*2048+ 836,   23*2048+1156,    0*2048+1601,
   0*2048+  99,    1*2048+1343,   33*2048+1387,    0*2048+1602,
   0*2048+ 111,   34*2048+ 188,   22*2048+ 869,    0*2048+1603,
   0*2048+ 122,   33*2048+ 123,   27*2048+ 541,    0*2048+1604,
   0*2048+ 132,   20*2048+ 254,   24*2048+1476,    0*2048+1605,
   0*2048+ 143,   29*2048+ 429,   17*2048+1299,    0*2048+1606,
   0*2048+ 155,   36*2048+ 265,   32*2048+1090,    0*2048+1607,
   0*2048+ 165,   27*2048+ 572,   23*2048+ 837,    0*2048+1608,
   0*2048+ 177,   35*2048+ 759,   31*2048+1013,    0*2048+1609,
  29*2048+  13,   34*2048+ 133,    0*2048+ 189,    0*2048+1610,
   0*2048+ 198,   15*2048+ 209,   18*2048+ 870,    0*2048+1620,
   0*2048+ 210,   10*2048+ 430,    9*2048+1122,    0*2048+1621,
   0*2048+ 221,   17*2048+ 794,   25*2048+1375,    0*2048+1622,
   0*2048+ 234,    7*2048+ 739,   27*2048+1111,    0*2048+1623,
   0*2048+ 243,   42*2048+ 352,   41*2048+1092,    0*2048+1624,
   0*2048+ 256,   12*2048+ 257,   41*2048+1565,    0*2048+1625,
   0*2048+ 266,   26*2048+ 662,   13*2048+ 903,    0*2048+1626,
   0*2048+ 277,    6*2048+1211,   29*2048+1477,    0*2048+1627,
   0*2048+ 288,   39*2048+1036,   23*2048+1355,    0*2048+1628,
  34*2048+   2,    0*2048+ 297,    1*2048+1543,    0*2048+1629,
   0*2048+ 309,   34*2048+ 386,   22*2048+1069,    0*2048+1630,
   0*2048+ 322,   33*2048+ 323,   27*2048+ 740,    0*2048+1631,
  25*2048+  91,    0*2048+ 330,   20*2048+ 452,    0*2048+1632,
   0*2048+ 342,   29*2048+ 628,   17*2048+1498,    0*2048+1633,
   0*2048+ 353,   36*2048+ 465,   32*2048+1290,    0*2048+1634,
   0*2048+ 363,   27*2048+ 771,   23*2048+1037,    0*2048+1635,
   0*2048+ 375,   35*2048+ 959,   31*2048+1212,    0*2048+1636,
  29*2048+ 211,   34*2048+ 331,    0*2048+ 387,    0*2048+1637,
   0*2048+ 396,   15*2048+ 409,   18*2048+1070,    0*2048+1647,
   0*2048+ 410,   10*2048+ 629,    9*2048+1321,    0*2048+1648,
   0*2048+ 421,   17*2048+ 993,   25*2048+1575,    0*2048+1649,
   0*2048+ 433,    7*2048+ 937,   27*2048+1309,    0*2048+1650,
   0*2048+ 441,   42*2048+ 550,   41*2048+1292,    0*2048+1651,
  42*2048+ 181,    0*2048+ 454,   12*2048+ 455,    0*2048+1652,
   0*2048+ 466,   26*2048+ 862,   13*2048+1102,    0*2048+1653,
  30*2048+  92,    0*2048+ 476,    6*2048+1411,    0*2048+1654,
   0*2048+ 487,   39*2048+1235,   23*2048+1554,    0*2048+1655,
   2*2048+ 159,   34*2048+ 200,    0*2048+ 495,    0*2048+1656,
   0*2048+ 508,   34*2048+ 585,   22*2048+1267,    0*2048+1657,
   0*2048+ 521,   33*2048+ 522,   27*2048+ 938,    0*2048+1658,
  25*2048+ 291,    0*2048+ 532,   20*2048+ 652,    0*2048+1659,
  18*2048+ 114,    0*2048+ 543,   29*2048+ 826,    0*2048+1660,
   0*2048+ 551,   36*2048+ 664,   32*2048+1489,    0*2048+1661,
   0*2048+ 562,   27*2048+ 969,   23*2048+1236,    0*2048+1662,
   0*2048+ 574,   35*2048+1159,   31*2048+1412,    0*2048+1663,
  29*2048+ 411,   34*2048+ 533,    0*2048+ 586,    0*2048+1664,
   0*2048+ 595,   15*2048+ 608,   18*2048+1268,    0*2048+1674,
   0*2048+ 609,   10*2048+ 827,    9*2048+1519,    0*2048+1675,
  26*2048+ 192,    0*2048+ 619,   17*2048+1193,    0*2048+1676,
   0*2048+ 632,    7*2048+1135,   27*2048+1509,    0*2048+1677,
   0*2048+ 640,   42*2048+ 750,   41*2048+1491,    0*2048+1678,
  42*2048+ 379,    0*2048+ 654,   12*2048+ 655,    0*2048+1679,
   0*2048+ 665,   26*2048+1060,   13*2048+1302,    0*2048+1680,
   7*2048+  26,   30*2048+ 292,    0*2048+ 675,    0*2048+1681,
  24*2048+ 169,    0*2048+ 686,   39*2048+1434,    0*2048+1682,
   2*2048+ 357,   34*2048+ 398,    0*2048+ 694,    0*2048+1683,
   0*2048+ 707,   34*2048+ 784,   22*2048+1466,    0*2048+1684,
   0*2048+ 719,   33*2048+ 720,   27*2048+1136,    0*2048+1685,
  25*2048+ 490,    0*2048+ 731,   20*2048+ 850,    0*2048+1686,
  18*2048+ 312,    0*2048+ 742,   29*2048+1024,    0*2048+1687,
  33*2048+ 104,    0*2048+ 751,   36*2048+ 864,    0*2048+1688,
   0*2048+ 761,   27*2048+1168,   23*2048+1435,    0*2048+1689,
  32*2048+  27,    0*2048+ 773,   35*2048+1358,    0*2048+1690,
  29*2048+ 610,   34*2048+ 732,    0*2048+ 785,    0*2048+1691,
   0*2048+ 795,   15*2048+ 807,   18*2048+1467,    0*2048+1701,
  10*2048+ 135,    0*2048+ 808,   10*2048+1025,    0*2048+1702,
  26*2048+ 390,    0*2048+ 817,   17*2048+1393,    0*2048+1703,
  28*2048+ 126,    0*2048+ 830,    7*2048+1335,    0*2048+1704,
  42*2048+ 106,    0*2048+ 840,   42*2048+ 948,    0*2048+1705,
  42*2048+ 578,    0*2048+ 852,   12*2048+ 853,    0*2048+1706,
   0*2048+ 865,   26*2048+1259,   13*2048+1501,    0*2048+1707,
   7*2048+ 225,   30*2048+ 491,    0*2048+ 874,    0*2048+1708,
  40*2048+  49,   24*2048+ 367,    0*2048+ 884,    0*2048+1709,
   2*2048+ 555,   34*2048+ 597,    0*2048+ 894,    0*2048+1710,
  23*2048+  82,    0*2048+ 906,   34*2048+ 983,    0*2048+1711,
   0*2048+ 918,   33*2048+ 919,   27*2048+1336,    0*2048+1712,
  25*2048+ 689,    0*2048+ 930,   20*2048+1048,    0*2048+1713,
  18*2048+ 511,    0*2048+ 940,   29*2048+1223,    0*2048+1714,
  33*2048+ 302,    0*2048+ 949,   36*2048+1062,    0*2048+1715,
  24*2048+  50,    0*2048+ 961,   27*2048+1369,    0*2048+1716,
  32*2048+ 226,    0*2048+ 971,   35*2048+1557,    0*2048+1717,
  29*2048+ 809,   34*2048+ 931,    0*2048+ 984,    0*2048+1718,
  19*2048+  83,    0*2048+ 994,   15*2048+1005,    0*2048+1728,
  10*2048+ 333,    0*2048+1006,   10*2048+1224,    0*2048+1729,
  18*2048+   8,   26*2048+ 589,    0*2048+1017,    0*2048+1730,
  28*2048+ 326,    0*2048+1028,    7*2048+1534,    0*2048+1731,
  42*2048+ 304,    0*2048+1040,   42*2048+1147,    0*2048+1732,
  42*2048+ 777,    0*2048+1050,   12*2048+1051,    0*2048+1733,
  14*2048+ 117,    0*2048+1063,   26*2048+1457,    0*2048+1734,
   7*2048+ 425,   30*2048+ 690,    0*2048+1074,    0*2048+1735,
  40*2048+ 248,   24*2048+ 566,    0*2048+1082,    0*2048+1736,
   2*2048+ 755,   34*2048+ 797,    0*2048+1094,    0*2048+1737,
  23*2048+ 281,    0*2048+1105,   34*2048+1182,    0*2048+1738,
   0*2048+1116,   33*2048+1117,   27*2048+1535,    0*2048+1739,
  25*2048+ 887,    0*2048+1128,   20*2048+1247,    0*2048+1740,
  18*2048+ 710,    0*2048+1138,   29*2048+1423,    0*2048+1741,
  33*2048+ 500,    0*2048+1148,   36*2048+1261,    0*2048+1742,
  24*2048+ 249,    0*2048+1161,   27*2048+1568,    0*2048+1743,
  36*2048+ 172,   32*2048+ 426,    0*2048+1170,    0*2048+1744,
  29*2048+1007,   34*2048+1129,    0*2048+1183,    0*2048+1745,
  19*2048+ 282,    0*2048+1194,   15*2048+1203,    0*2048+1755,
  10*2048+ 535,    0*2048+1204,   10*2048+1424,    0*2048+1756,
  18*2048+ 206,   26*2048+ 788,    0*2048+1216,    0*2048+1757,
   8*2048+ 149,   28*2048+ 525,    0*2048+1227,    0*2048+1758,
  42*2048+ 502,    0*2048+1239,   42*2048+1347,    0*2048+1759,
  42*2048+ 975,    0*2048+1249,   12*2048+1250,    0*2048+1760,
  27*2048+  72,   14*2048+ 315,    0*2048+1262,    0*2048+1761,
   7*2048+ 623,   30*2048+ 888,    0*2048+1272,    0*2048+1762,
  40*2048+ 446,   24*2048+ 765,    0*2048+1281,    0*2048+1763,
   2*2048+ 953,   34*2048+ 996,    0*2048+1294,    0*2048+1764,
  23*2048+ 480,    0*2048+1305,   34*2048+1380,    0*2048+1765,
  28*2048+ 150,    0*2048+1314,   33*2048+1315,    0*2048+1766,
  25*2048+1085,    0*2048+1327,   20*2048+1446,    0*2048+1767,
  30*2048+  40,   18*2048+ 909,    0*2048+1338,    0*2048+1768,
  33*2048+ 699,    0*2048+1348,   36*2048+1459,    0*2048+1769,
  28*2048+ 184,   24*2048+ 447,    0*2048+1360,    0*2048+1770,
  36*2048+ 370,   32*2048+ 624,    0*2048+1371,    0*2048+1771,
  29*2048+1205,   34*2048+1328,    0*2048+1381,    0*2048+1772,
  19*2048+ 481,    0*2048+1394,   15*2048+1403,    0*2048+1782,
  11*2048+  41,   10*2048+ 734,    0*2048+1404,    0*2048+1783,
  18*2048+ 404,   26*2048+ 987,    0*2048+1416,    0*2048+1784,
   8*2048+ 348,   28*2048+ 723,    0*2048+1427,    0*2048+1785,
  42*2048+ 701,    0*2048+1438,   42*2048+1547,    0*2048+1786,
  42*2048+1174,    0*2048+1448,   12*2048+1449,    0*2048+1787,
  27*2048+ 272,   14*2048+ 514,    0*2048+1460,    0*2048+1788,
   7*2048+ 821,   30*2048+1086,    0*2048+1471,    0*2048+1789,
  40*2048+ 645,   24*2048+ 965,    0*2048+1482,    0*2048+1790,
   2*2048+1152,   34*2048+1196,    0*2048+1493,    0*2048+1791,
  23*2048+ 679,    0*2048+1504,   34*2048+1580,    0*2048+1792,
  28*2048+ 349,    0*2048+1514,   33*2048+1515,    0*2048+1793,
  21*2048+  63,   25*2048+1284,    0*2048+1525,    0*2048+1794,
  30*2048+ 239,   18*2048+1108,    0*2048+1537,    0*2048+1795,
  37*2048+  74,   33*2048+ 899,    0*2048+1548,    0*2048+1796,
  28*2048+ 382,   24*2048+ 646,    0*2048+1559,    0*2048+1797,
  36*2048+ 569,   32*2048+ 822,    0*2048+1570,    0*2048+1798,
  29*2048+1405,   34*2048+1526,    0*2048+1581,    0*2048+1799,
  15*2048+ 242,   19*2048+ 319,    5*2048+ 561,   33*2048+ 649,    9*2048+ 858,   23*2048+ 902,   44*2048+ 990,   39*2048+1067,   19*2048+1144,    3*2048+1232,   29*2048+1474,   24*2048+1540,    0*2048+1584,
   5*2048+  33,   18*2048+ 253,   15*2048+ 528,   20*2048+ 529,   34*2048+ 605,    1*2048+ 737,   41*2048+ 979,    8*2048+1034,    2*2048+1210,    1*2048+1331,   39*2048+1353,   38*2048+1419,    0*2048+1585,
  40*2048+ 187,   34*2048+ 473,   43*2048+ 506,    1*2048+ 726,   21*2048+ 792,   29*2048+1166,    7*2048+1221,   36*2048+1254,   32*2048+1342,   44*2048+1397,   43*2048+1408,   27*2048+1409,    0*2048+1586,
  33*2048+  55,   14*2048+ 517,   39*2048+ 530,   27*2048+ 748,   23*2048+1100,   29*2048+1188,    3*2048+1441,   21*2048+1463,   28*2048+1485,   16*2048+1507,   41*2048+1551,   43*2048+1562,    0*2048+1587,
  43*2048+  34,   31*2048+ 110,    5*2048+ 176,   29*2048+ 275,    0*2048+ 650,   26*2048+ 693,   10*2048+ 803,   20*2048+1287,   16*2048+1364,   32*2048+1365,   11*2048+1508,    2*2048+1541,    0*2048+1588,
  30*2048+ 462,   44*2048+ 531,   40*2048+ 539,   21*2048+ 627,   26*2048+ 682,   31*2048+ 770,   18*2048+ 859,   37*2048+ 891,   35*2048+1089,   13*2048+1398,   40*2048+1420,   25*2048+1496,    0*2048+1589,
  16*2048+  77,    6*2048+ 121,   20*2048+ 286,   40*2048+ 407,   11*2048+ 418,   38*2048+ 484,    8*2048+ 583,   26*2048+ 793,   24*2048+ 957,    5*2048+1068,    8*2048+1155,   22*2048+1288,    0*2048+1590,
  15*2048+ 264,   39*2048+ 287,   16*2048+ 320,   29*2048+ 749,   37*2048+ 958,    7*2048+1243,   41*2048+1298,   12*2048+1320,   11*2048+1332,   33*2048+1475,   24*2048+1529,    1*2048+1573,    0*2048+1591,
   6*2048+ 220,   27*2048+ 341,   28*2048+ 408,   39*2048+ 419,   12*2048+ 638,    9*2048+ 660,   20*2048+ 781,   19*2048+1035,    2*2048+1189,   14*2048+1386,   32*2048+1430,    8*2048+1574,    0*2048+1592,
  30*2048+  89,   25*2048+ 156,   15*2048+ 440,   19*2048+ 518,    5*2048+ 760,   33*2048+ 847,    9*2048+1056,   23*2048+1101,   44*2048+1190,   39*2048+1265,   19*2048+1344,    3*2048+1431,    0*2048+1611,
  39*2048+  36,    5*2048+ 232,   18*2048+ 451,   15*2048+ 727,   20*2048+ 728,   34*2048+ 804,    1*2048+ 935,   41*2048+1178,    8*2048+1233,    2*2048+1410,    1*2048+1530,   39*2048+1552,    0*2048+1612,
  45*2048+  14,   44*2048+  23,   28*2048+  24,   40*2048+ 385,   34*2048+ 672,   43*2048+ 705,    1*2048+ 925,   21*2048+ 991,   29*2048+1367,    7*2048+1421,   36*2048+1452,   32*2048+1542,    0*2048+1613,
   4*2048+  58,   22*2048+  79,   29*2048+ 100,   17*2048+ 124,   42*2048+ 166,   44*2048+ 178,   33*2048+ 255,   14*2048+ 715,   39*2048+ 729,   27*2048+ 946,   23*2048+1300,   29*2048+1388,    0*2048+1614,
  12*2048+ 125,    3*2048+ 157,   43*2048+ 233,   31*2048+ 308,    5*2048+ 374,   29*2048+ 474,    0*2048+ 848,   26*2048+ 893,   10*2048+1001,   20*2048+1486,   16*2048+1563,   32*2048+1564,    0*2048+1615,
  14*2048+  15,   41*2048+  37,   26*2048+ 112,   30*2048+ 661,   44*2048+ 730,   40*2048+ 738,   21*2048+ 825,   26*2048+ 880,   31*2048+ 968,   18*2048+1057,   37*2048+1091,   35*2048+1289,    0*2048+1616,
  16*2048+ 276,    6*2048+ 321,   20*2048+ 485,   40*2048+ 606,   11*2048+ 616,   38*2048+ 683,    8*2048+ 782,   26*2048+ 992,   24*2048+1157,    5*2048+1266,    8*2048+1354,   22*2048+1487,    0*2048+1617,
  34*2048+  90,   25*2048+ 144,    2*2048+ 190,   15*2048+ 464,   39*2048+ 486,   16*2048+ 519,   29*2048+ 947,   37*2048+1158,    7*2048+1442,   41*2048+1497,   12*2048+1518,   11*2048+1531,    0*2048+1618,
  15*2048+   1,   33*2048+  45,    9*2048+ 191,    6*2048+ 420,   27*2048+ 542,   28*2048+ 607,   39*2048+ 617,   12*2048+ 838,    9*2048+ 860,   20*2048+ 980,   19*2048+1234,    2*2048+1389,    0*2048+1619,
   4*2048+  46,   30*2048+ 289,   25*2048+ 354,   15*2048+ 639,   19*2048+ 716,    5*2048+ 960,   33*2048+1045,    9*2048+1255,   23*2048+1301,   44*2048+1390,   39*2048+1464,   19*2048+1544,    0*2048+1638,
   3*2048+  25,    2*2048+ 145,   40*2048+ 167,   39*2048+ 235,    5*2048+ 431,   18*2048+ 651,   15*2048+ 926,   20*2048+ 927,   34*2048+1002,    1*2048+1133,   41*2048+1376,    8*2048+1432,    0*2048+1639,
   8*2048+  38,   37*2048+  67,   33*2048+ 158,   45*2048+ 212,   44*2048+ 222,   28*2048+ 223,   40*2048+ 584,   34*2048+ 871,   43*2048+ 904,    1*2048+1123,   21*2048+1191,   29*2048+1566,    0*2048+1640,
  30*2048+   3,    4*2048+ 258,   22*2048+ 278,   29*2048+ 298,   17*2048+ 324,   42*2048+ 364,   44*2048+ 376,   33*2048+ 453,   14*2048+ 914,   39*2048+ 928,   27*2048+1145,   23*2048+1499,    0*2048+1641,
  21*2048+ 101,   17*2048+ 179,   33*2048+ 180,   12*2048+ 325,    3*2048+ 355,   43*2048+ 432,   31*2048+ 507,    5*2048+ 573,   29*2048+ 673,    0*2048+1046,   26*2048+1093,   10*2048+1199,    0*2048+1642,
  14*2048+ 213,   41*2048+ 236,   26*2048+ 310,   30*2048+ 861,   44*2048+ 929,   40*2048+ 936,   21*2048+1023,   26*2048+1078,   31*2048+1167,   18*2048+1256,   37*2048+1291,   35*2048+1488,    0*2048+1643,
  23*2048+ 102,   16*2048+ 475,    6*2048+ 520,   20*2048+ 684,   40*2048+ 805,   11*2048+ 814,   38*2048+ 881,    8*2048+ 981,   26*2048+1192,   24*2048+1356,    5*2048+1465,    8*2048+1553,    0*2048+1644,
   8*2048+  59,   42*2048+ 113,   13*2048+ 134,   12*2048+ 146,   34*2048+ 290,   25*2048+ 343,    2*2048+ 388,   15*2048+ 663,   39*2048+ 685,   16*2048+ 717,   29*2048+1146,   37*2048+1357,    0*2048+1645,
   3*2048+   4,   15*2048+ 199,   33*2048+ 244,    9*2048+ 389,    6*2048+ 618,   27*2048+ 741,   28*2048+ 806,   39*2048+ 815,   12*2048+1038,    9*2048+1058,   20*2048+1179,   19*2048+1433,    0*2048+1646,
  45*2048+   5,   40*2048+  80,   20*2048+ 160,    4*2048+ 245,   30*2048+ 488,   25*2048+ 552,   15*2048+ 839,   19*2048+ 915,    5*2048+1160,   33*2048+1244,    9*2048+1453,   23*2048+1500,    0*2048+1665,
   9*2048+  47,    3*2048+ 224,    2*2048+ 344,   40*2048+ 365,   39*2048+ 434,    5*2048+ 630,   18*2048+ 849,   15*2048+1124,   20*2048+1125,   34*2048+1200,    1*2048+1333,   41*2048+1576,    0*2048+1666,
  30*2048+ 182,    8*2048+ 237,   37*2048+ 267,   33*2048+ 356,   45*2048+ 412,   44*2048+ 422,   28*2048+ 423,   40*2048+ 783,   34*2048+1071,   43*2048+1103,    1*2048+1322,   21*2048+1391,    0*2048+1667,
  24*2048+ 115,   30*2048+ 201,    4*2048+ 456,   22*2048+ 477,   29*2048+ 496,   17*2048+ 523,   42*2048+ 563,   44*2048+ 575,   33*2048+ 653,   14*2048+1112,   39*2048+1126,   27*2048+1345,    0*2048+1668,
  21*2048+ 299,   17*2048+ 377,   33*2048+ 378,   12*2048+ 524,    3*2048+ 553,   43*2048+ 631,   31*2048+ 706,    5*2048+ 772,   29*2048+ 872,    0*2048+1245,   26*2048+1293,   10*2048+1399,    0*2048+1669,
  36*2048+ 103,   14*2048+ 413,   41*2048+ 435,   26*2048+ 509,   30*2048+1059,   44*2048+1127,   40*2048+1134,   21*2048+1222,   26*2048+1277,   31*2048+1368,   18*2048+1454,   37*2048+1490,    0*2048+1670,
   6*2048+  81,    9*2048+ 168,   23*2048+ 300,   16*2048+ 674,    6*2048+ 718,   20*2048+ 882,   40*2048+1003,   11*2048+1014,   38*2048+1079,    8*2048+1180,   26*2048+1392,   24*2048+1555,    0*2048+1671,
   8*2048+ 259,   42*2048+ 311,   13*2048+ 332,   12*2048+ 345,   34*2048+ 489,   25*2048+ 544,    2*2048+ 587,   15*2048+ 863,   39*2048+ 883,   16*2048+ 916,   29*2048+1346,   37*2048+1556,    0*2048+1672,
  20*2048+  48,    3*2048+ 202,   15*2048+ 397,   33*2048+ 442,    9*2048+ 588,    6*2048+ 816,   27*2048+ 939,   28*2048+1004,   39*2048+1015,   12*2048+1237,    9*2048+1257,   20*2048+1377,    0*2048+1673,
  10*2048+  68,   24*2048+ 116,   45*2048+ 203,   40*2048+ 279,   20*2048+ 358,    4*2048+ 443,   30*2048+ 687,   25*2048+ 752,   15*2048+1039,   19*2048+1113,    5*2048+1359,   33*2048+1443,    0*2048+1692,
  42*2048+ 193,    9*2048+ 246,    3*2048+ 424,    2*2048+ 545,   40*2048+ 564,   39*2048+ 633,    5*2048+ 828,   18*2048+1047,   15*2048+1323,   20*2048+1324,   34*2048+1400,    1*2048+1532,    0*2048+1693,
  22*2048+   6,   30*2048+ 380,    8*2048+ 436,   37*2048+ 467,   33*2048+ 554,   45*2048+ 611,   44*2048+ 620,   28*2048+ 621,   40*2048+ 982,   34*2048+1269,   43*2048+1303,    1*2048+1520,    0*2048+1694,
  24*2048+ 313,   30*2048+ 399,    4*2048+ 656,   22*2048+ 676,   29*2048+ 695,   17*2048+ 721,   42*2048+ 762,   44*2048+ 774,   33*2048+ 851,   14*2048+1310,   39*2048+1325,   27*2048+1545,    0*2048+1695,
  11*2048+  16,   21*2048+ 497,   17*2048+ 576,   33*2048+ 577,   12*2048+ 722,    3*2048+ 753,   43*2048+ 829,   31*2048+ 905,    5*2048+ 970,   29*2048+1072,    0*2048+1444,   26*2048+1492,    0*2048+1696,
  19*2048+  69,   38*2048+ 105,   36*2048+ 301,   14*2048+ 612,   41*2048+ 634,   26*2048+ 708,   30*2048+1258,   44*2048+1326,   40*2048+1334,   21*2048+1422,   26*2048+1478,   31*2048+1567,    0*2048+1697,
  27*2048+   7,   25*2048+ 170,    6*2048+ 280,    9*2048+ 366,   23*2048+ 498,   16*2048+ 873,    6*2048+ 917,   20*2048+1080,   40*2048+1201,   11*2048+1213,   38*2048+1278,    8*2048+1378,    0*2048+1698,
  38*2048+ 171,    8*2048+ 457,   42*2048+ 510,   13*2048+ 534,   12*2048+ 546,   34*2048+ 688,   25*2048+ 743,    2*2048+ 786,   15*2048+1061,   39*2048+1081,   16*2048+1114,   29*2048+1546,    0*2048+1699,
  20*2048+ 247,    3*2048+ 400,   15*2048+ 596,   33*2048+ 641,    9*2048+ 787,    6*2048+1016,   27*2048+1137,   28*2048+1202,   39*2048+1214,   12*2048+1436,    9*2048+1455,   20*2048+1577,    0*2048+1700,
  34*2048+  60,   10*2048+ 268,   24*2048+ 314,   45*2048+ 401,   40*2048+ 478,   20*2048+ 556,    4*2048+ 642,   30*2048+ 885,   25*2048+ 950,   15*2048+1238,   19*2048+1311,    5*2048+1558,    0*2048+1719,
  35*2048+  17,    2*2048+ 147,   42*2048+ 391,    9*2048+ 444,    3*2048+ 622,    2*2048+ 744,   40*2048+ 763,   39*2048+ 831,    5*2048+1026,   18*2048+1246,   15*2048+1521,   20*2048+1522,    0*2048+1720,
   2*2048+ 136,   22*2048+ 204,   30*2048+ 579,    8*2048+ 635,   37*2048+ 666,   33*2048+ 754,   45*2048+ 810,   44*2048+ 818,   28*2048+ 819,   40*2048+1181,   34*2048+1468,   43*2048+1502,    0*2048+1721,
  28*2048+ 161,   24*2048+ 512,   30*2048+ 598,    4*2048+ 854,   22*2048+ 875,   29*2048+ 895,   17*2048+ 920,   42*2048+ 962,   44*2048+ 972,   33*2048+1049,   14*2048+1510,   39*2048+1523,    0*2048+1722,
   1*2048+  61,   27*2048+ 107,   11*2048+ 214,   21*2048+ 696,   17*2048+ 775,   33*2048+ 776,   12*2048+ 921,    3*2048+ 951,   43*2048+1027,   31*2048+1104,    5*2048+1169,   29*2048+1270,    0*2048+1723,
  22*2048+  39,   27*2048+  93,   32*2048+ 183,   19*2048+ 269,   38*2048+ 303,   36*2048+ 499,   14*2048+ 811,   41*2048+ 832,   26*2048+ 907,   30*2048+1456,   44*2048+1524,   40*2048+1533,    0*2048+1724,
  27*2048+ 205,   25*2048+ 368,    6*2048+ 479,    9*2048+ 565,   23*2048+ 697,   16*2048+1073,    6*2048+1115,   20*2048+1279,   40*2048+1401,   11*2048+1413,   38*2048+1479,    8*2048+1578,    0*2048+1725,
  30*2048+ 162,   38*2048+ 369,    8*2048+ 657,   42*2048+ 709,   13*2048+ 733,   12*2048+ 745,   34*2048+ 886,   25*2048+ 941,    2*2048+ 985,   15*2048+1260,   39*2048+1280,   16*2048+1312,    0*2048+1726,
  13*2048+  51,   10*2048+  70,   21*2048+ 194,   20*2048+ 445,    3*2048+ 599,   15*2048+ 796,   33*2048+ 841,    9*2048+ 986,    6*2048+1215,   27*2048+1337,   28*2048+1402,   39*2048+1414,    0*2048+1727,
   6*2048+ 173,   34*2048+ 260,   10*2048+ 468,   24*2048+ 513,   45*2048+ 600,   40*2048+ 677,   20*2048+ 756,    4*2048+ 842,   30*2048+1083,   25*2048+1149,   15*2048+1437,   19*2048+1511,    0*2048+1746,
  16*2048+ 137,   21*2048+ 138,   35*2048+ 215,    2*2048+ 346,   42*2048+ 590,    9*2048+ 643,    3*2048+ 820,    2*2048+ 942,   40*2048+ 963,   39*2048+1029,    5*2048+1225,   18*2048+1445,    0*2048+1747,
  35*2048+  84,   44*2048+ 118,    2*2048+ 334,   22*2048+ 402,   30*2048+ 778,    8*2048+ 833,   37*2048+ 866,   33*2048+ 952,   45*2048+1008,   44*2048+1018,   28*2048+1019,   40*2048+1379,    0*2048+1748,
  15*2048+ 127,   40*2048+ 139,   28*2048+ 359,   24*2048+ 711,   30*2048+ 798,    4*2048+1052,   22*2048+1075,   29*2048+1095,   17*2048+1118,   42*2048+1162,   44*2048+1171,   33*2048+1248,    0*2048+1749,
   1*2048+ 261,   27*2048+ 305,   11*2048+ 414,   21*2048+ 896,   17*2048+ 973,   33*2048+ 974,   12*2048+1119,    3*2048+1150,   43*2048+1226,   31*2048+1304,    5*2048+1370,   29*2048+1469,    0*2048+1750,
  31*2048+  71,   45*2048+ 140,   41*2048+ 148,   22*2048+ 238,   27*2048+ 293,   32*2048+ 381,   19*2048+ 469,   38*2048+ 501,   36*2048+ 698,   14*2048+1009,   41*2048+1030,   26*2048+1106,    0*2048+1751,
  41*2048+  18,   12*2048+  28,   39*2048+  94,    9*2048+ 195,   27*2048+ 403,   25*2048+ 567,    6*2048+ 678,    9*2048+ 764,   23*2048+ 897,   16*2048+1271,    6*2048+1313,   20*2048+1480,    0*2048+1752,
  30*2048+ 360,   38*2048+ 568,    8*2048+ 855,   42*2048+ 908,   13*2048+ 932,   12*2048+ 943,   34*2048+1084,   25*2048+1139,    2*2048+1184,   15*2048+1458,   39*2048+1481,   16*2048+1512,    0*2048+1753,
  29*2048+  19,   40*2048+  29,   13*2048+ 250,   10*2048+ 270,   21*2048+ 392,   20*2048+ 644,    3*2048+ 799,   15*2048+ 995,   33*2048+1041,    9*2048+1185,    6*2048+1415,   27*2048+1536,    0*2048+1754,
  16*2048+  52,   20*2048+ 128,    6*2048+ 371,   34*2048+ 458,   10*2048+ 667,   24*2048+ 712,   45*2048+ 800,   40*2048+ 876,   20*2048+ 954,    4*2048+1042,   30*2048+1282,   25*2048+1349,    0*2048+1773,
  19*2048+  62,   16*2048+ 335,   21*2048+ 336,   35*2048+ 415,    2*2048+ 547,   42*2048+ 789,    9*2048+ 843,    3*2048+1020,    2*2048+1140,   40*2048+1163,   39*2048+1228,    5*2048+1425,    0*2048+1774,
  35*2048+ 283,   44*2048+ 316,    2*2048+ 536,   22*2048+ 601,   30*2048+ 976,    8*2048+1031,   37*2048+1064,   33*2048+1151,   45*2048+1206,   44*2048+1217,   28*2048+1218,   40*2048+1579,    0*2048+1775,
  15*2048+ 327,   40*2048+ 337,   28*2048+ 557,   24*2048+ 910,   30*2048+ 997,    4*2048+1251,   22*2048+1273,   29*2048+1295,   17*2048+1316,   42*2048+1361,   44*2048+1372,   33*2048+1447,    0*2048+1776,
  30*2048+  85,    1*2048+ 459,   27*2048+ 503,   11*2048+ 613,   21*2048+1096,   17*2048+1172,   33*2048+1173,   12*2048+1317,    3*2048+1350,   43*2048+1426,   31*2048+1503,    5*2048+1569,    0*2048+1777,
  31*2048+ 271,   45*2048+ 338,   41*2048+ 347,   22*2048+ 437,   27*2048+ 492,   32*2048+ 580,   19*2048+ 668,   38*2048+ 700,   36*2048+ 898,   14*2048+1207,   41*2048+1229,   26*2048+1306,    0*2048+1778,
  21*2048+  95,   41*2048+ 216,   12*2048+ 227,   39*2048+ 294,    9*2048+ 393,   27*2048+ 602,   25*2048+ 766,    6*2048+ 877,    9*2048+ 964,   23*2048+1097,   16*2048+1470,    6*2048+1513,    0*2048+1779,
  16*2048+  73,   40*2048+  96,   17*2048+ 129,   30*2048+ 558,   38*2048+ 767,    8*2048+1053,   42*2048+1107,   13*2048+1130,   12*2048+1141,   34*2048+1283,   25*2048+1339,    2*2048+1382,    0*2048+1780,
   7*2048+  30,   28*2048+ 151,   29*2048+ 217,   40*2048+ 228,   13*2048+ 448,   10*2048+ 470,   21*2048+ 591,   20*2048+ 844,    3*2048+ 998,   15*2048+1195,   33*2048+1240,    9*2048+1383,    0*2048+1781,

   0*2048+   8,    0*2048+  18,    0*2048+1440,
   0*2048+  19,    0*2048+  28,    0*2048+1441,
   0*2048+  29,    0*2048+  38,    0*2048+1442,
   0*2048+  39,    0*2048+  48,    0*2048+1443,
   0*2048+  49,    0*2048+  58,    0*2048+1444,
   0*2048+  59,    0*2048+  68,    0*2048+1445,
   0*2048+  69,    0*2048+  78,    0*2048+1446,
   0*2048+  79,    0*2048+  88,    0*2048+1447,
   0*2048+  89,    0*2048+  98,    0*2048+1448,
   0*2048+  99,    0*2048+ 108,    0*2048+1449,
   0*2048+ 109,    0*2048+ 118,    0*2048+1450,
   0*2048+ 119,    0*2048+ 128,    0*2048+1451,
   0*2048+ 129,    0*2048+ 138,    0*2048+1452,
   0*2048+ 139,    0*2048+ 148,    0*2048+1453,
   0*2048+ 149,    0*2048+ 158,    0*2048+1454,
   0*2048+ 159,    0*2048+ 168,    0*2048+1455,
   0*2048+ 169,    0*2048+ 178,    0*2048+1456,
   0*2048+ 179,    0*2048+ 188,    0*2048+1457,
   0*2048+ 189,    0*2048+ 198,    0*2048+1458,
   0*2048+ 199,    0*2048+ 208,    0*2048+1459,
   0*2048+ 209,    0*2048+ 218,    0*2048+1460,
   0*2048+ 219,    0*2048+ 228,    0*2048+1461,
   0*2048+ 229,    0*2048+ 238,    0*2048+1462,
   0*2048+ 239,    0*2048+ 248,    0*2048+1463,
   0*2048+ 249,    0*2048+ 258,    0*2048+1464,
   0*2048+ 259,    0*2048+ 268,    0*2048+1465,
   0*2048+ 269,    0*2048+ 278,    0*2048+1466,
   0*2048+ 279,    0*2048+ 288,    0*2048+1467,
   0*2048+ 289,    0*2048+ 298,    0*2048+1468,
   0*2048+ 299,    0*2048+ 308,    0*2048+1469,
   0*2048+ 309,    0*2048+ 318,    0*2048+1470,
   0*2048+ 319,    0*2048+ 328,    0*2048+1471,
   0*2048+ 329,    0*2048+ 338,    0*2048+1472,
   0*2048+ 339,    0*2048+ 348,    0*2048+1473,
   0*2048+ 349,    0*2048+ 358,    0*2048+1474,
   0*2048+ 359,    0*2048+ 368,    0*2048+1475,
   0*2048+ 369,    0*2048+ 378,    0*2048+1476,
   0*2048+ 379,    0*2048+ 388,    0*2048+1477,
   0*2048+ 389,    0*2048+ 398,    0*2048+1478,
   0*2048+ 399,    0*2048+ 408,    0*2048+1479,
   0*2048+ 409,    0*2048+ 418,    0*2048+1480,
   0*2048+ 419,    0*2048+ 428,    0*2048+1481,
   0*2048+ 429,    0*2048+ 438,    0*2048+1482,
   0*2048+ 439,    0*2048+ 448,    0*2048+1483,
   0*2048+ 449,    0*2048+ 458,    0*2048+1484,
   0*2048+ 459,    0*2048+ 468,    0*2048+1485,
   0*2048+ 469,    0*2048+ 478,    0*2048+1486,
   0*2048+ 479,    0*2048+ 488,    0*2048+1487,
   0*2048+ 489,    0*2048+ 498,    0*2048+1488,
   0*2048+ 499,    0*2048+ 508,    0*2048+1489,
   0*2048+ 509,    0*2048+ 518,    0*2048+1490,
   0*2048+ 519,    0*2048+ 528,    0*2048+1491,
   0*2048+ 529,    0*2048+ 538,    0*2048+1492,
   0*2048+ 539,    0*2048+ 548,    0*2048+1493,
   0*2048+ 549,    0*2048+ 558,    0*2048+1494,
   0*2048+ 559,    0*2048+ 568,    0*2048+1495,
   0*2048+ 569,    0*2048+ 578,    0*2048+1496,
   0*2048+ 579,    0*2048+ 588,    0*2048+1497,
   0*2048+ 589,    0*2048+ 598,    0*2048+1498,
   0*2048+ 599,    0*2048+ 608,    0*2048+1499,
   0*2048+ 609,    0*2048+ 618,    0*2048+1500,
   0*2048+ 619,    0*2048+ 628,    0*2048+1501,
   0*2048+ 629,    0*2048+ 638,    0*2048+1502,
   0*2048+ 639,    0*2048+ 648,    0*2048+1503,
   0*2048+ 649,    0*2048+ 658,    0*2048+1504,
   0*2048+ 659,    0*2048+ 668,    0*2048+1505,
   0*2048+ 669,    0*2048+ 678,    0*2048+1506,
   0*2048+ 679,    0*2048+ 688,    0*2048+1507,
   0*2048+ 689,    0*2048+ 698,    0*2048+1508,
   0*2048+ 699,    0*2048+ 708,    0*2048+1509,
   0*2048+ 709,    0*2048+ 718,    0*2048+1510,
   0*2048+ 719,    0*2048+ 728,    0*2048+1511,
   0*2048+ 729,    0*2048+ 738,    0*2048+1512,
   0*2048+ 739,    0*2048+ 748,    0*2048+1513,
   0*2048+ 749,    0*2048+ 758,    0*2048+1514,
   0*2048+ 759,    0*2048+ 768,    0*2048+1515,
   0*2048+ 769,    0*2048+ 778,    0*2048+1516,
   0*2048+ 779,    0*2048+ 788,    0*2048+1517,
   0*2048+ 789,    0*2048+ 798,    0*2048+1518,
   0*2048+ 799,    0*2048+ 808,    0*2048+1519,
   0*2048+ 809,    0*2048+ 818,    0*2048+1520,
   0*2048+ 819,    0*2048+ 828,    0*2048+1521,
   0*2048+ 829,    0*2048+ 838,    0*2048+1522,
   0*2048+ 839,    0*2048+ 848,    0*2048+1523,
   0*2048+ 849,    0*2048+ 858,    0*2048+1524,
   0*2048+ 859,    0*2048+ 868,    0*2048+1525,
   0*2048+ 869,    0*2048+ 878,    0*2048+1526,
   0*2048+ 879,    0*2048+ 888,    0*2048+1527,
   0*2048+ 889,    0*2048+ 898,    0*2048+1528,
   0*2048+ 899,    0*2048+ 908,    0*2048+1529,
   0*2048+ 909,    0*2048+ 918,    0*2048+1530,
   0*2048+ 919,    0*2048+ 928,    0*2048+1531,
   0*2048+ 929,    0*2048+ 938,    0*2048+1532,
   0*2048+ 939,    0*2048+ 948,    0*2048+1533,
   0*2048+ 949,    0*2048+ 958,    0*2048+1534,
   0*2048+ 959,    0*2048+ 968,    0*2048+1535,
   0*2048+ 969,    0*2048+ 978,    0*2048+1536,
   0*2048+ 979,    0*2048+ 988,    0*2048+1537,
   0*2048+ 989,    0*2048+ 998,    0*2048+1538,
   0*2048+ 999,    0*2048+1008,    0*2048+1539,
   0*2048+1009,    0*2048+1018,    0*2048+1540,
   0*2048+1019,    0*2048+1028,    0*2048+1541,
   0*2048+1029,    0*2048+1038,    0*2048+1542,
   0*2048+1039,    0*2048+1048,    0*2048+1543,
   0*2048+1049,    0*2048+1058,    0*2048+1544,
   0*2048+1059,    0*2048+1068,    0*2048+1545,
   0*2048+1069,    0*2048+1078,    0*2048+1546,
   0*2048+1079,    0*2048+1088,    0*2048+1547,
   0*2048+1089,    0*2048+1098,    0*2048+1548,
   0*2048+1099,    0*2048+1108,    0*2048+1549,
   0*2048+1109,    0*2048+1118,    0*2048+1550,
   0*2048+1119,    0*2048+1128,    0*2048+1551,
   0*2048+1129,    0*2048+1138,    0*2048+1552,
   0*2048+1139,    0*2048+1148,    0*2048+1553,
   0*2048+1149,    0*2048+1158,    0*2048+1554,
   0*2048+1159,    0*2048+1168,    0*2048+1555,
   0*2048+1169,    0*2048+1178,    0*2048+1556,
   0*2048+1179,    0*2048+1188,    0*2048+1557,
   0*2048+1189,    0*2048+1198,    0*2048+1558,
   1*2048+   9,    0*2048+1199,    0*2048+1559,
   0*2048+  30,   29*2048+ 491,    2*2048+1021,    0*2048+1203,
   0*2048+  40,   17*2048+1071,   34*2048+1180,    0*2048+1204,
   0*2048+  51,   40*2048+ 361,   15*2048+ 800,    0*2048+1205,
   0*2048+  60,   32*2048+ 241,   40*2048+1100,    0*2048+1206,
   2*2048+  31,    0*2048+  71,   12*2048+1022,    0*2048+1207,
   0*2048+  80,   25*2048+ 111,   11*2048+1160,    0*2048+1208,
  18*2048+  72,    0*2048+  91,   20*2048+1120,    0*2048+1209,
   0*2048+ 101,    8*2048+ 430,   38*2048+ 460,    0*2048+1210,
   0*2048+ 112,   23*2048+ 750,    5*2048+1050,    0*2048+1211,
   0*2048+ 120,   28*2048+ 660,   19*2048+ 850,    0*2048+1212,
  32*2048+  81,    0*2048+ 131,   20*2048+ 740,    0*2048+1213,
   0*2048+ 140,   11*2048+ 400,   14*2048+ 630,    0*2048+1214,
   0*2048+   2,   21*2048+ 160,    1*2048+ 431,    0*2048+1215,
   0*2048+  11,   21*2048+ 631,    9*2048+1000,    0*2048+1216,
   0*2048+  22,    4*2048+ 290,   12*2048+1023,    0*2048+1217,
   0*2048+  32,    8*2048+ 450,   36*2048+ 980,    0*2048+1218,
   0*2048+  41,   43*2048+ 520,   42*2048+ 770,    0*2048+1219,
   0*2048+  52,   24*2048+ 420,   17*2048+1150,    0*2048+1220,
   0*2048+  61,   22*2048+ 560,    2*2048+1072,    0*2048+1221,
   0*2048+  73,   35*2048+ 960,    1*2048+1060,    0*2048+1222,
  13*2048+   3,    4*2048+  74,    0*2048+  82,    0*2048+1223,
   0*2048+  92,   13*2048+ 801,   32*2048+ 861,    0*2048+1224,
   0*2048+ 102,    1*2048+ 291,   24*2048+ 480,    0*2048+1225,
   0*2048+ 113,    4*2048+ 830,   19*2048+ 840,    0*2048+1226,
   0*2048+ 121,    5*2048+ 350,    5*2048+ 881,    0*2048+1227,
  14*2048+  42,    0*2048+ 132,    1*2048+1110,    0*2048+1228,
   0*2048+ 141,    9*2048+ 492,   32*2048+ 540,    0*2048+1229,
   0*2048+ 180,   29*2048+ 641,    2*2048+1171,    0*2048+1233,
  18*2048+  24,   35*2048+ 133,    0*2048+ 191,    0*2048+1234,
   0*2048+ 202,   40*2048+ 511,   15*2048+ 950,    0*2048+1235,
  41*2048+  53,    0*2048+ 210,   32*2048+ 392,    0*2048+1236,
   2*2048+ 181,    0*2048+ 221,   12*2048+1172,    0*2048+1237,
  12*2048+ 114,    0*2048+ 230,   25*2048+ 261,    0*2048+1238,
  21*2048+  75,   18*2048+ 222,    0*2048+ 243,    0*2048+1239,
   0*2048+ 251,    8*2048+ 580,   38*2048+ 610,    0*2048+1240,
   6*2048+   4,    0*2048+ 262,   23*2048+ 900,    0*2048+1241,
   0*2048+ 270,   28*2048+ 811,   19*2048+1001,    0*2048+1242,
  32*2048+ 231,    0*2048+ 281,   20*2048+ 891,    0*2048+1243,
   0*2048+ 292,   11*2048+ 550,   14*2048+ 780,    0*2048+1244,
   0*2048+ 152,   21*2048+ 310,    1*2048+ 581,    0*2048+1245,
   0*2048+ 162,   21*2048+ 781,    9*2048+1151,    0*2048+1246,
   0*2048+ 172,    4*2048+ 442,   12*2048+1173,    0*2048+1247,
   0*2048+ 182,    8*2048+ 601,   36*2048+1131,    0*2048+1248,
   0*2048+ 192,   43*2048+ 670,   42*2048+ 920,    0*2048+1249,
  18*2048+ 103,    0*2048+ 203,   24*2048+ 570,    0*2048+1250,
   3*2048+  25,    0*2048+ 211,   22*2048+ 710,    0*2048+1251,
   2*2048+  12,    0*2048+ 223,   35*2048+1111,    0*2048+1252,
  13*2048+ 153,    4*2048+ 224,    0*2048+ 232,    0*2048+1253,
   0*2048+ 244,   13*2048+ 951,   32*2048+1011,    0*2048+1254,
   0*2048+ 252,    1*2048+ 443,   24*2048+ 632,    0*2048+1255,
   0*2048+ 263,    4*2048+ 981,   19*2048+ 990,    0*2048+1256,
   0*2048+ 271,    5*2048+ 500,    5*2048+1031,    0*2048+1257,
   2*2048+  62,   14*2048+ 193,    0*2048+ 282,    0*2048+1258,
   0*2048+ 293,    9*2048+ 642,   32*2048+ 690,    0*2048+1259,
   3*2048+ 123,    0*2048+ 330,   29*2048+ 792,    0*2048+1263,
  18*2048+ 174,   35*2048+ 283,    0*2048+ 341,    0*2048+1264,
   0*2048+ 353,   40*2048+ 662,   15*2048+1101,    0*2048+1265,
  41*2048+ 204,    0*2048+ 362,   32*2048+ 543,    0*2048+1266,
  13*2048+ 124,    2*2048+ 331,    0*2048+ 371,    0*2048+1267,
  12*2048+ 264,    0*2048+ 381,   25*2048+ 411,    0*2048+1268,
  21*2048+ 225,   18*2048+ 372,    0*2048+ 394,    0*2048+1269,
   0*2048+ 402,    8*2048+ 730,   38*2048+ 762,    0*2048+1270,
   6*2048+ 154,    0*2048+ 412,   23*2048+1051,    0*2048+1271,
   0*2048+ 421,   28*2048+ 962,   19*2048+1152,    0*2048+1272,
  32*2048+ 382,    0*2048+ 433,   20*2048+1041,    0*2048+1273,
   0*2048+ 444,   11*2048+ 701,   14*2048+ 930,    0*2048+1274,
   0*2048+ 302,   21*2048+ 461,    1*2048+ 731,    0*2048+1275,
  10*2048+ 104,    0*2048+ 312,   21*2048+ 931,    0*2048+1276,
  13*2048+ 125,    0*2048+ 322,    4*2048+ 592,    0*2048+1277,
  37*2048+  84,    0*2048+ 332,    8*2048+ 752,    0*2048+1278,
   0*2048+ 342,   43*2048+ 820,   42*2048+1073,    0*2048+1279,
  18*2048+ 253,    0*2048+ 354,   24*2048+ 720,    0*2048+1280,
   3*2048+ 175,    0*2048+ 363,   22*2048+ 862,    0*2048+1281,
  36*2048+  63,    2*2048+ 163,    0*2048+ 373,    0*2048+1282,
  13*2048+ 303,    4*2048+ 374,    0*2048+ 383,    0*2048+1283,
   0*2048+ 395,   13*2048+1102,   32*2048+1162,    0*2048+1284,
   0*2048+ 403,    1*2048+ 593,   24*2048+ 782,    0*2048+1285,
   0*2048+ 413,    4*2048+1132,   19*2048+1140,    0*2048+1286,
   0*2048+ 422,    5*2048+ 650,    5*2048+1182,    0*2048+1287,
   2*2048+ 212,   14*2048+ 343,    0*2048+ 434,    0*2048+1288,
   0*2048+ 445,    9*2048+ 793,   32*2048+ 841,    0*2048+1289,
   3*2048+ 273,    0*2048+ 481,   29*2048+ 942,    0*2048+1293,
  18*2048+ 324,   35*2048+ 435,    0*2048+ 494,    0*2048+1294,
  16*2048+  54,    0*2048+ 503,   40*2048+ 813,    0*2048+1295,
  41*2048+ 355,    0*2048+ 512,   32*2048+ 693,    0*2048+1296,
  13*2048+ 274,    2*2048+ 482,    0*2048+ 522,    0*2048+1297,
  12*2048+ 414,    0*2048+ 532,   25*2048+ 562,    0*2048+1298,
  21*2048+ 375,   18*2048+ 523,    0*2048+ 545,    0*2048+1299,
   0*2048+ 552,    8*2048+ 882,   38*2048+ 913,    0*2048+1300,
  24*2048+   5,    6*2048+ 304,    0*2048+ 563,    0*2048+1301,
  20*2048+ 105,    0*2048+ 571,   28*2048+1113,    0*2048+1302,
  32*2048+ 533,    0*2048+ 583,   20*2048+1191,    0*2048+1303,
   0*2048+ 594,   11*2048+ 852,   14*2048+1082,    0*2048+1304,
   0*2048+ 453,   21*2048+ 611,    1*2048+ 883,    0*2048+1305,
  10*2048+ 254,    0*2048+ 463,   21*2048+1083,    0*2048+1306,
  13*2048+ 275,    0*2048+ 473,    4*2048+ 743,    0*2048+1307,
  37*2048+ 234,    0*2048+ 483,    8*2048+ 902,    0*2048+1308,
  43*2048+  26,    0*2048+ 495,   43*2048+ 971,    0*2048+1309,
  18*2048+ 404,    0*2048+ 504,   24*2048+ 871,    0*2048+1310,
   3*2048+ 325,    0*2048+ 513,   22*2048+1012,    0*2048+1311,
  36*2048+ 213,    2*2048+ 313,    0*2048+ 524,    0*2048+1312,
  13*2048+ 454,    4*2048+ 525,    0*2048+ 534,    0*2048+1313,
  14*2048+  55,   33*2048+ 116,    0*2048+ 546,    0*2048+1314,
   0*2048+ 553,    1*2048+ 744,   24*2048+ 932,    0*2048+1315,
   5*2048+  85,   20*2048+  93,    0*2048+ 564,    0*2048+1316,
   6*2048+ 135,    0*2048+ 572,    5*2048+ 802,    0*2048+1317,
   2*2048+ 364,   14*2048+ 496,    0*2048+ 584,    0*2048+1318,
   0*2048+ 595,    9*2048+ 943,   32*2048+ 991,    0*2048+1319,
   3*2048+ 424,    0*2048+ 633,   29*2048+1092,    0*2048+1323,
  18*2048+ 475,   35*2048+ 585,    0*2048+ 644,    0*2048+1324,
  16*2048+ 205,    0*2048+ 653,   40*2048+ 964,    0*2048+1325,
  41*2048+ 505,    0*2048+ 663,   32*2048+ 844,    0*2048+1326,
  13*2048+ 425,    2*2048+ 634,    0*2048+ 672,    0*2048+1327,
  12*2048+ 565,    0*2048+ 682,   25*2048+ 712,    0*2048+1328,
  21*2048+ 526,   18*2048+ 673,    0*2048+ 695,    0*2048+1329,
   0*2048+ 703,    8*2048+1032,   38*2048+1064,    0*2048+1330,
  24*2048+ 155,    6*2048+ 455,    0*2048+ 713,    0*2048+1331,
  29*2048+  65,   20*2048+ 255,    0*2048+ 721,    0*2048+1332,
  21*2048+ 143,   32*2048+ 683,    0*2048+ 733,    0*2048+1333,
  15*2048+  35,    0*2048+ 745,   11*2048+1003,    0*2048+1334,
   0*2048+ 604,   21*2048+ 763,    1*2048+1033,    0*2048+1335,
  22*2048+  36,   10*2048+ 405,    0*2048+ 613,    0*2048+1336,
  13*2048+ 426,    0*2048+ 623,    4*2048+ 894,    0*2048+1337,
  37*2048+ 385,    0*2048+ 635,    8*2048+1053,    0*2048+1338,
  43*2048+ 176,    0*2048+ 645,   43*2048+1122,    0*2048+1339,
  18*2048+ 554,    0*2048+ 654,   24*2048+1025,    0*2048+1340,
   3*2048+ 476,    0*2048+ 664,   22*2048+1163,    0*2048+1341,
  36*2048+ 365,    2*2048+ 464,    0*2048+ 674,    0*2048+1342,
  13*2048+ 605,    4*2048+ 675,    0*2048+ 684,    0*2048+1343,
  14*2048+ 206,   33*2048+ 266,    0*2048+ 696,    0*2048+1344,
   0*2048+ 704,    1*2048+ 895,   24*2048+1084,    0*2048+1345,
   5*2048+ 235,   20*2048+ 245,    0*2048+ 714,    0*2048+1346,
   6*2048+ 285,    0*2048+ 722,    5*2048+ 952,    0*2048+1347,
   2*2048+ 514,   14*2048+ 646,    0*2048+ 734,    0*2048+1348,
   0*2048+ 746,    9*2048+1093,   32*2048+1141,    0*2048+1349,
  30*2048+  45,    3*2048+ 574,    0*2048+ 783,    0*2048+1353,
  18*2048+ 625,   35*2048+ 735,    0*2048+ 795,    0*2048+1354,
  16*2048+ 356,    0*2048+ 805,   40*2048+1115,    0*2048+1355,
  41*2048+ 655,    0*2048+ 814,   32*2048+ 994,    0*2048+1356,
  13*2048+ 575,    2*2048+ 784,    0*2048+ 822,    0*2048+1357,
  12*2048+ 715,    0*2048+ 833,   25*2048+ 864,    0*2048+1358,
  21*2048+ 676,   18*2048+ 823,    0*2048+ 846,    0*2048+1359,
  39*2048+  16,    0*2048+ 854,    8*2048+1183,    0*2048+1360,
  24*2048+ 305,    6*2048+ 606,    0*2048+ 865,    0*2048+1361,
  29*2048+ 215,   20*2048+ 406,    0*2048+ 872,    0*2048+1362,
  21*2048+ 295,   32*2048+ 834,    0*2048+ 885,    0*2048+1363,
  15*2048+ 185,    0*2048+ 896,   11*2048+1154,    0*2048+1364,
   0*2048+ 755,   21*2048+ 914,    1*2048+1184,    0*2048+1365,
  22*2048+ 186,   10*2048+ 555,    0*2048+ 765,    0*2048+1366,
  13*2048+ 576,    0*2048+ 774,    4*2048+1044,    0*2048+1367,
   9*2048+   7,   37*2048+ 536,    0*2048+ 785,    0*2048+1368,
  44*2048+  77,   43*2048+ 326,    0*2048+ 796,    0*2048+1369,
  18*2048+ 705,    0*2048+ 806,   24*2048+1175,    0*2048+1370,
  23*2048+ 117,    3*2048+ 626,    0*2048+ 815,    0*2048+1371,
  36*2048+ 515,    2*2048+ 614,    0*2048+ 824,    0*2048+1372,
  13*2048+ 756,    4*2048+ 825,    0*2048+ 835,    0*2048+1373,
  14*2048+ 357,   33*2048+ 416,    0*2048+ 847,    0*2048+1374,
  25*2048+  37,    0*2048+ 855,    1*2048+1045,    0*2048+1375,
   5*2048+ 386,   20*2048+ 396,    0*2048+ 866,    0*2048+1376,
   6*2048+ 437,    0*2048+ 873,    5*2048+1103,    0*2048+1377,
   2*2048+ 665,   14*2048+ 797,    0*2048+ 886,    0*2048+1378,
  10*2048+  46,   33*2048+  94,    0*2048+ 897,    0*2048+1379,
  30*2048+ 196,    3*2048+ 724,    0*2048+ 933,    0*2048+1383,
  18*2048+ 776,   35*2048+ 887,    0*2048+ 945,    0*2048+1384,
  41*2048+  67,   16*2048+ 506,    0*2048+ 955,    0*2048+1385,
  41*2048+ 807,    0*2048+ 965,   32*2048+1144,    0*2048+1386,
  13*2048+ 725,    2*2048+ 934,    0*2048+ 973,    0*2048+1387,
  12*2048+ 867,    0*2048+ 984,   25*2048+1014,    0*2048+1388,
  21*2048+ 826,   18*2048+ 974,    0*2048+ 996,    0*2048+1389,
   9*2048+ 136,   39*2048+ 167,    0*2048+1005,    0*2048+1390,
  24*2048+ 456,    6*2048+ 757,    0*2048+1015,    0*2048+1391,
  29*2048+ 367,   20*2048+ 556,    0*2048+1026,    0*2048+1392,
  21*2048+ 447,   32*2048+ 985,    0*2048+1035,    0*2048+1393,
  12*2048+ 107,   15*2048+ 335,    0*2048+1046,    0*2048+1394,
   2*2048+ 137,    0*2048+ 905,   21*2048+1065,    0*2048+1395,
  22*2048+ 336,   10*2048+ 706,    0*2048+ 916,    0*2048+1396,
  13*2048+ 726,    0*2048+ 924,    4*2048+1194,    0*2048+1397,
   9*2048+ 157,   37*2048+ 686,    0*2048+ 935,    0*2048+1398,
  44*2048+ 227,   43*2048+ 477,    0*2048+ 946,    0*2048+1399,
  25*2048+ 127,   18*2048+ 856,    0*2048+ 956,    0*2048+1400,
  23*2048+ 267,    3*2048+ 777,    0*2048+ 966,    0*2048+1401,
  36*2048+ 666,    2*2048+ 766,    0*2048+ 975,    0*2048+1402,
  13*2048+ 906,    4*2048+ 976,    0*2048+ 986,    0*2048+1403,
  14*2048+ 507,   33*2048+ 567,    0*2048+ 997,    0*2048+1404,
  25*2048+ 187,    0*2048+1006,    1*2048+1195,    0*2048+1405,
   5*2048+ 537,   20*2048+ 547,    0*2048+1016,    0*2048+1406,
   6*2048+  56,    6*2048+ 587,    0*2048+1027,    0*2048+1407,
   2*2048+ 816,   14*2048+ 947,    0*2048+1036,    0*2048+1408,
  10*2048+ 197,   33*2048+ 246,    0*2048+1047,    0*2048+1409,
  30*2048+ 346,    3*2048+ 875,    0*2048+1085,    0*2048+1413,
  18*2048+ 926,   35*2048+1037,    0*2048+1095,    0*2048+1414,
  41*2048+ 217,   16*2048+ 656,    0*2048+1106,    0*2048+1415,
  33*2048+  97,   41*2048+ 957,    0*2048+1116,    0*2048+1416,
  13*2048+ 876,    2*2048+1086,    0*2048+1124,    0*2048+1417,
  12*2048+1017,    0*2048+1135,   25*2048+1165,    0*2048+1418,
  21*2048+ 977,   18*2048+1125,    0*2048+1146,    0*2048+1419,
   9*2048+ 286,   39*2048+ 317,    0*2048+1156,    0*2048+1420,
  24*2048+ 607,    6*2048+ 907,    0*2048+1166,    0*2048+1421,
  29*2048+ 517,   20*2048+ 707,    0*2048+1176,    0*2048+1422,
  21*2048+ 597,   32*2048+1136,    0*2048+1186,    0*2048+1423,
  12*2048+ 257,   15*2048+ 486,    0*2048+1196,    0*2048+1424,
  22*2048+  17,    2*2048+ 287,    0*2048+1056,    0*2048+1425,
  22*2048+ 487,   10*2048+ 857,    0*2048+1067,    0*2048+1426,
   5*2048+ 146,   13*2048+ 877,    0*2048+1077,    0*2048+1427,
   9*2048+ 307,   37*2048+ 837,    0*2048+1087,    0*2048+1428,
  44*2048+ 377,   43*2048+ 627,    0*2048+1096,    0*2048+1429,
  25*2048+ 277,   18*2048+1007,    0*2048+1107,    0*2048+1430,
  23*2048+ 417,    3*2048+ 927,    0*2048+1117,    0*2048+1431,
  36*2048+ 817,    2*2048+ 917,    0*2048+1126,    0*2048+1432,
  13*2048+1057,    4*2048+1127,    0*2048+1137,    0*2048+1433,
  14*2048+ 657,   33*2048+ 717,    0*2048+1147,    0*2048+1434,
   2*2048+ 147,   25*2048+ 337,    0*2048+1157,    0*2048+1435,
   5*2048+ 687,   20*2048+ 697,    0*2048+1167,    0*2048+1436,
   6*2048+ 207,    6*2048+ 737,    0*2048+1177,    0*2048+1437,
   2*2048+ 967,   14*2048+1097,    0*2048+1187,    0*2048+1438,
  10*2048+ 347,   33*2048+ 397,    0*2048+1197,    0*2048+1439,
   0*2048+   0,   28*2048+  90,   12*2048+ 200,   17*2048+ 440,   13*2048+ 530,   38*2048+ 600,   26*2048+ 760,   20*2048+ 810,   10*2048+ 860,   28*2048+ 910,   35*2048+ 970,   21*2048+1020,   12*2048+1080,    0*2048+1200,
  24*2048+   1,    0*2048+  10,    1*2048+  20,    8*2048+ 110,    3*2048+ 130,   36*2048+ 380,   15*2048+ 470,   29*2048+ 490,   12*2048+ 761,   31*2048+ 790,   11*2048+ 870,   28*2048+ 880,   25*2048+1081,    0*2048+1201,
   0*2048+  21,   26*2048+  50,   44*2048+  70,   22*2048+ 100,    2*2048+ 190,    7*2048+ 240,   33*2048+ 360,   28*2048+ 390,    1*2048+ 441,   19*2048+ 700,    7*2048+ 890,    0*2048+1070,   31*2048+1130,    0*2048+1202,
  13*2048+  33,    0*2048+ 150,   28*2048+ 242,   12*2048+ 351,   17*2048+ 590,   13*2048+ 680,   38*2048+ 751,   26*2048+ 911,   20*2048+ 961,   10*2048+1010,   28*2048+1061,   35*2048+1121,   21*2048+1170,    0*2048+1230,
  26*2048+  34,   24*2048+ 151,    0*2048+ 161,    1*2048+ 170,    8*2048+ 260,    3*2048+ 280,   36*2048+ 531,   15*2048+ 620,   29*2048+ 640,   12*2048+ 912,   31*2048+ 940,   11*2048+1024,   28*2048+1030,    0*2048+1231,
   1*2048+  23,   32*2048+  83,    0*2048+ 171,   26*2048+ 201,   44*2048+ 220,   22*2048+ 250,    2*2048+ 340,    7*2048+ 391,   33*2048+ 510,   28*2048+ 541,    1*2048+ 591,   19*2048+ 851,    7*2048+1040,    0*2048+1232,
  29*2048+  13,   36*2048+  76,   22*2048+ 122,   13*2048+ 183,    0*2048+ 300,   28*2048+ 393,   12*2048+ 501,   17*2048+ 741,   13*2048+ 831,   38*2048+ 901,   26*2048+1062,   20*2048+1112,   10*2048+1161,    0*2048+1260,
  26*2048+ 184,   24*2048+ 301,    0*2048+ 311,    1*2048+ 320,    8*2048+ 410,    3*2048+ 432,   36*2048+ 681,   15*2048+ 771,   29*2048+ 791,   12*2048+1063,   31*2048+1090,   11*2048+1174,   28*2048+1181,    0*2048+1261,
   1*2048+ 173,   32*2048+ 233,    0*2048+ 321,   26*2048+ 352,   44*2048+ 370,   22*2048+ 401,    2*2048+ 493,    7*2048+ 542,   33*2048+ 661,   28*2048+ 691,    1*2048+ 742,   19*2048+1002,    7*2048+1190,    0*2048+1262,
  27*2048+  14,   21*2048+  64,   11*2048+ 115,   29*2048+ 164,   36*2048+ 226,   22*2048+ 272,   13*2048+ 333,    0*2048+ 451,   28*2048+ 544,   12*2048+ 651,   17*2048+ 892,   13*2048+ 982,   38*2048+1052,    0*2048+1290,
  13*2048+  15,   32*2048+  43,   12*2048+ 126,   29*2048+ 134,   26*2048+ 334,   24*2048+ 452,    0*2048+ 462,    1*2048+ 471,    8*2048+ 561,    3*2048+ 582,   36*2048+ 832,   15*2048+ 921,   29*2048+ 941,    0*2048+1291,
   8*2048+ 142,    1*2048+ 323,   32*2048+ 384,    0*2048+ 472,   26*2048+ 502,   44*2048+ 521,   22*2048+ 551,    2*2048+ 643,    7*2048+ 692,   33*2048+ 812,   28*2048+ 842,    1*2048+ 893,   19*2048+1153,    0*2048+1292,
  39*2048+   6,   27*2048+ 165,   21*2048+ 214,   11*2048+ 265,   29*2048+ 314,   36*2048+ 376,   22*2048+ 423,   13*2048+ 484,    0*2048+ 602,   28*2048+ 694,   12*2048+ 803,   17*2048+1042,   13*2048+1133,    0*2048+1320,
  13*2048+ 166,   32*2048+ 194,   12*2048+ 276,   29*2048+ 284,   26*2048+ 485,   24*2048+ 603,    0*2048+ 612,    1*2048+ 621,    8*2048+ 711,    3*2048+ 732,   36*2048+ 983,   15*2048+1074,   29*2048+1091,    0*2048+1321,
  20*2048+ 106,    8*2048+ 294,    1*2048+ 474,   32*2048+ 535,    0*2048+ 622,   26*2048+ 652,   44*2048+ 671,   22*2048+ 702,    2*2048+ 794,    7*2048+ 843,   33*2048+ 963,   28*2048+ 992,    1*2048+1043,    0*2048+1322,
  14*2048+  86,   39*2048+ 156,   27*2048+ 315,   21*2048+ 366,   11*2048+ 415,   29*2048+ 465,   36*2048+ 527,   22*2048+ 573,   13*2048+ 636,    0*2048+ 753,   28*2048+ 845,   12*2048+ 953,   17*2048+1192,    0*2048+1350,
  16*2048+  27,   30*2048+  44,   13*2048+ 316,   32*2048+ 344,   12*2048+ 427,   29*2048+ 436,   26*2048+ 637,   24*2048+ 754,    0*2048+ 764,    1*2048+ 772,    8*2048+ 863,    3*2048+ 884,   36*2048+1134,    0*2048+1351,
  20*2048+ 256,    8*2048+ 446,    1*2048+ 624,   32*2048+ 685,    0*2048+ 773,   26*2048+ 804,   44*2048+ 821,   22*2048+ 853,    2*2048+ 944,    7*2048+ 993,   33*2048+1114,   28*2048+1142,    1*2048+1193,    0*2048+1352,
  18*2048+ 144,   14*2048+ 236,   39*2048+ 306,   27*2048+ 466,   21*2048+ 516,   11*2048+ 566,   29*2048+ 615,   36*2048+ 677,   22*2048+ 723,   13*2048+ 786,    0*2048+ 903,   28*2048+ 995,   12*2048+1104,    0*2048+1380,
  37*2048+  87,   16*2048+ 177,   30*2048+ 195,   13*2048+ 467,   32*2048+ 497,   12*2048+ 577,   29*2048+ 586,   26*2048+ 787,   24*2048+ 904,    0*2048+ 915,    1*2048+ 922,    8*2048+1013,    3*2048+1034,    0*2048+1381,
  34*2048+  66,   29*2048+  95,    2*2048+ 145,   20*2048+ 407,    8*2048+ 596,    1*2048+ 775,   32*2048+ 836,    0*2048+ 923,   26*2048+ 954,   44*2048+ 972,   22*2048+1004,    2*2048+1094,    7*2048+1143,    0*2048+1382,
  13*2048+  57,   18*2048+ 296,   14*2048+ 387,   39*2048+ 457,   27*2048+ 616,   21*2048+ 667,   11*2048+ 716,   29*2048+ 767,   36*2048+ 827,   22*2048+ 874,   13*2048+ 936,    0*2048+1054,   28*2048+1145,    0*2048+1410,
  37*2048+ 237,   16*2048+ 327,   30*2048+ 345,   13*2048+ 617,   32*2048+ 647,   12*2048+ 727,   29*2048+ 736,   26*2048+ 937,   24*2048+1055,    0*2048+1066,    1*2048+1075,    8*2048+1164,    3*2048+1185,    0*2048+1411,
   3*2048+  47,    8*2048+  96,   34*2048+ 216,   29*2048+ 247,    2*2048+ 297,   20*2048+ 557,    8*2048+ 747,    1*2048+ 925,   32*2048+ 987,    0*2048+1076,   26*2048+1105,   44*2048+1123,   22*2048+1155,    0*2048+1412,

   0*2048+   8,    0*2048+  20,    0*2048+1320,
   0*2048+  21,    0*2048+  31,    0*2048+1321,
   0*2048+  32,    0*2048+  40,    0*2048+1322,
   0*2048+  41,    0*2048+  50,    0*2048+1323,
   0*2048+  51,    0*2048+  63,    0*2048+1324,
   0*2048+  64,    0*2048+  74,    0*2048+1325,
   0*2048+  75,    0*2048+  86,    0*2048+1326,
   0*2048+  87,    0*2048+  97,    0*2048+1327,
   0*2048+  98,    0*2048+ 107,    0*2048+1328,
   0*2048+ 108,    0*2048+ 118,    0*2048+1329,
   0*2048+ 119,    0*2048+ 130,    0*2048+1330,
   0*2048+ 131,    0*2048+ 140,    0*2048+1331,
   0*2048+ 141,    0*2048+ 152,    0*2048+1332,
   0*2048+ 153,    0*2048+ 163,    0*2048+1333,
   0*2048+ 164,    0*2048+ 172,    0*2048+1334,
   0*2048+ 173,    0*2048+ 182,    0*2048+1335,
   0*2048+ 183,    0*2048+ 195,    0*2048+1336,
   0*2048+ 196,    0*2048+ 206,    0*2048+1337,
   0*2048+ 207,    0*2048+ 218,    0*2048+1338,
   0*2048+ 219,    0*2048+ 229,    0*2048+1339,
   0*2048+ 230,    0*2048+ 239,    0*2048+1340,
   0*2048+ 240,    0*2048+ 250,    0*2048+1341,
   0*2048+ 251,    0*2048+ 262,    0*2048+1342,
   0*2048+ 263,    0*2048+ 272,    0*2048+1343,
   0*2048+ 273,    0*2048+ 284,    0*2048+1344,
   0*2048+ 285,    0*2048+ 295,    0*2048+1345,
   0*2048+ 296,    0*2048+ 304,    0*2048+1346,
   0*2048+ 305,    0*2048+ 314,    0*2048+1347,
   0*2048+ 315,    0*2048+ 327,    0*2048+1348,
   0*2048+ 328,    0*2048+ 338,    0*2048+1349,
   0*2048+ 339,    0*2048+ 350,    0*2048+1350,
   0*2048+ 351,    0*2048+ 361,    0*2048+1351,
   0*2048+ 362,    0*2048+ 371,    0*2048+1352,
   0*2048+ 372,    0*2048+ 382,    0*2048+1353,
   0*2048+ 383,    0*2048+ 394,    0*2048+1354,
   0*2048+ 395,    0*2048+ 404,    0*2048+1355,
   0*2048+ 405,    0*2048+ 416,    0*2048+1356,
   0*2048+ 417,    0*2048+ 427,    0*2048+1357,
   0*2048+ 428,    0*2048+ 436,    0*2048+1358,
   0*2048+ 437,    0*2048+ 446,    0*2048+1359,
   0*2048+ 447,    0*2048+ 459,    0*2048+1360,
   0*2048+ 460,    0*2048+ 470,    0*2048+1361,
   0*2048+ 471,    0*2048+ 482,    0*2048+1362,
   0*2048+ 483,    0*2048+ 493,    0*2048+1363,
   0*2048+ 494,    0*2048+ 503,    0*2048+1364,
   0*2048+ 504,    0*2048+ 514,    0*2048+1365,
   0*2048+ 515,    0*2048+ 526,    0*2048+1366,
   0*2048+ 527,    0*2048+ 536,    0*2048+1367,
   0*2048+ 537,    0*2048+ 548,    0*2048+1368,
   0*2048+ 549,    0*2048+ 559,    0*2048+1369,
   0*2048+ 560,    0*2048+ 568,    0*2048+1370,
   0*2048+ 569,    0*2048+ 578,    0*2048+1371,
   0*2048+ 579,    0*2048+ 591,    0*2048+1372,
   0*2048+ 592,    0*2048+ 602,    0*2048+1373,
   0*2048+ 603,    0*2048+ 614,    0*2048+1374,
   0*2048+ 615,    0*2048+ 625,    0*2048+1375,
   0*2048+ 626,    0*2048+ 635,    0*2048+1376,
   0*2048+ 636,    0*2048+ 646,    0*2048+1377,
   0*2048+ 647,    0*2048+ 658,    0*2048+1378,
   0*2048+ 659,    0*2048+ 668,    0*2048+1379,
   0*2048+ 669,    0*2048+ 680,    0*2048+1380,
   0*2048+ 681,    0*2048+ 691,    0*2048+1381,
   0*2048+ 692,    0*2048+ 700,    0*2048+1382,
   0*2048+ 701,    0*2048+ 710,    0*2048+1383,
   0*2048+ 711,    0*2048+ 723,    0*2048+1384,
   0*2048+ 724,    0*2048+ 734,    0*2048+1385,
   0*2048+ 735,    0*2048+ 746,    0*2048+1386,
   0*2048+ 747,    0*2048+ 757,    0*2048+1387,
   0*2048+ 758,    0*2048+ 767,    0*2048+1388,
   0*2048+ 768,    0*2048+ 778,    0*2048+1389,
   0*2048+ 779,    0*2048+ 790,    0*2048+1390,
   0*2048+ 791,    0*2048+ 800,    0*2048+1391,
   0*2048+ 801,    0*2048+ 812,    0*2048+1392,
   0*2048+ 813,    0*2048+ 823,    0*2048+1393,
   0*2048+ 824,    0*2048+ 832,    0*2048+1394,
   0*2048+ 833,    0*2048+ 842,    0*2048+1395,
   0*2048+ 843,    0*2048+ 855,    0*2048+1396,
   0*2048+ 856,    0*2048+ 866,    0*2048+1397,
   0*2048+ 867,    0*2048+ 878,    0*2048+1398,
   0*2048+ 879,    0*2048+ 889,    0*2048+1399,
   0*2048+ 890,    0*2048+ 899,    0*2048+1400,
   0*2048+ 900,    0*2048+ 910,    0*2048+1401,
   0*2048+ 911,    0*2048+ 922,    0*2048+1402,
   0*2048+ 923,    0*2048+ 932,    0*2048+1403,
   0*2048+ 933,    0*2048+ 944,    0*2048+1404,
   0*2048+ 945,    0*2048+ 955,    0*2048+1405,
   0*2048+ 956,    0*2048+ 964,    0*2048+1406,
   0*2048+ 965,    0*2048+ 974,    0*2048+1407,
   0*2048+ 975,    0*2048+ 987,    0*2048+1408,
   0*2048+ 988,    0*2048+ 998,    0*2048+1409,
   0*2048+ 999,    0*2048+1010,    0*2048+1410,
   0*2048+1011,    0*2048+1021,    0*2048+1411,
   0*2048+1022,    0*2048+1031,    0*2048+1412,
   0*2048+1032,    0*2048+1042,    0*2048+1413,
   0*2048+1043,    0*2048+1054,    0*2048+1414,
   1*2048+   9,    0*2048+1055,    0*2048+1415,
   0*2048+  43,   22*2048+ 252,   27*2048+ 976,    0*2048+1057,
   0*2048+  52,   32*2048+ 384,   41*2048+1000,    0*2048+1058,
   0*2048+  65,   35*2048+ 142,   27*2048+ 495,    0*2048+1059,
   0*2048+  76,   39*2048+ 946,   35*2048+ 977,    0*2048+1060,
  43*2048+  10,    0*2048+  88,   21*2048+ 484,    0*2048+1061,
   0*2048+  99,   28*2048+ 593,   43*2048+ 616,    0*2048+1062,
   0*2048+ 109,   41*2048+ 110,   11*2048+ 154,    0*2048+1063,
   0*2048+ 121,   10*2048+ 265,   23*2048+ 340,    0*2048+1064,
   0*2048+   0,   15*2048+ 197,   31*2048+ 604,    0*2048+1065,
   0*2048+  11,   31*2048+ 297,   13*2048+ 880,    0*2048+1066,
   0*2048+  22,   11*2048+ 891,   17*2048+ 924,    0*2048+1067,
   0*2048+  34,    1*2048+ 396,   38*2048+ 845,    0*2048+1068,
   0*2048+  44,    6*2048+ 682,   18*2048+ 978,    0*2048+1069,
   0*2048+  53,   18*2048+ 505,   35*2048+ 957,    0*2048+1070,
   0*2048+  66,   13*2048+ 100,   37*2048+ 881,    0*2048+1071,
   0*2048+  77,   38*2048+ 506,    5*2048+ 683,    0*2048+1072,
   0*2048+  89,   20*2048+ 274,   10*2048+ 605,    0*2048+1073,
   0*2048+ 101,   20*2048+ 306,    4*2048+ 307,    0*2048+1074,
   0*2048+ 111,   23*2048+ 330,   10*2048+ 385,    0*2048+1075,
   0*2048+ 122,   43*2048+ 143,   19*2048+ 912,    0*2048+1076,
   0*2048+   1,   32*2048+  78,   25*2048+ 882,    0*2048+1077,
   0*2048+  12,   11*2048+ 352,   31*2048+ 496,    0*2048+1078,
   0*2048+  23,   14*2048+ 386,    7*2048+ 449,    0*2048+1079,
   0*2048+  35,   10*2048+ 406,   40*2048+ 693,    0*2048+1080,
  35*2048+  13,    0*2048+  45,   24*2048+ 208,    0*2048+1081,
   0*2048+  54,   10*2048+ 286,   11*2048+ 594,    0*2048+1082,
   0*2048+  67,   26*2048+ 397,    1*2048+ 507,    0*2048+1083,
  25*2048+  55,    0*2048+  79,   17*2048+ 637,    0*2048+1084,
   0*2048+  90,   13*2048+ 550,   19*2048+ 627,    0*2048+1085,
   0*2048+ 102,    6*2048+ 429,    1*2048+ 857,    0*2048+1086,
   0*2048+ 112,   17*2048+ 174,   32*2048+ 438,    0*2048+1087,
   0*2048+ 123,   29*2048+ 266,   14*2048+ 780,    0*2048+1088,
  28*2048+  56,    0*2048+ 176,   22*2048+ 387,    0*2048+1090,
  42*2048+  80,    0*2048+ 184,   32*2048+ 516,    0*2048+1091,
   0*2048+ 198,   35*2048+ 275,   27*2048+ 628,    0*2048+1092,
  40*2048+  24,   36*2048+  57,    0*2048+ 209,    0*2048+1093,
  43*2048+ 144,    0*2048+ 220,   21*2048+ 617,    0*2048+1094,
   0*2048+ 231,   28*2048+ 725,   43*2048+ 748,    0*2048+1095,
   0*2048+ 241,   41*2048+ 242,   11*2048+ 287,    0*2048+1096,
   0*2048+ 254,   10*2048+ 399,   23*2048+ 472,    0*2048+1097,
   0*2048+ 132,   15*2048+ 331,   31*2048+ 736,    0*2048+1098,
   0*2048+ 145,   31*2048+ 430,   13*2048+1012,    0*2048+1099,
  18*2048+   2,    0*2048+ 155,   11*2048+1023,    0*2048+1100,
   0*2048+ 166,    1*2048+ 528,   38*2048+ 980,    0*2048+1101,
  19*2048+  58,    0*2048+ 177,    6*2048+ 815,    0*2048+1102,
  36*2048+  36,    0*2048+ 185,   18*2048+ 638,    0*2048+1103,
   0*2048+ 199,   13*2048+ 232,   37*2048+1013,    0*2048+1104,
   0*2048+ 210,   38*2048+ 639,    5*2048+ 816,    0*2048+1105,
   0*2048+ 221,   20*2048+ 407,   10*2048+ 737,    0*2048+1106,
   0*2048+ 233,   20*2048+ 439,    4*2048+ 440,    0*2048+1107,
   0*2048+ 243,   23*2048+ 462,   10*2048+ 517,    0*2048+1108,
   0*2048+ 255,   43*2048+ 276,   19*2048+1044,    0*2048+1109,
   0*2048+ 133,   32*2048+ 211,   25*2048+1014,    0*2048+1110,
   0*2048+ 146,   11*2048+ 485,   31*2048+ 629,    0*2048+1111,
   0*2048+ 156,   14*2048+ 518,    7*2048+ 581,    0*2048+1112,
   0*2048+ 167,   10*2048+ 539,   40*2048+ 825,    0*2048+1113,
  35*2048+ 147,    0*2048+ 178,   24*2048+ 341,    0*2048+1114,
   0*2048+ 186,   10*2048+ 418,   11*2048+ 726,    0*2048+1115,
   0*2048+ 200,   26*2048+ 529,    1*2048+ 640,    0*2048+1116,
  25*2048+ 187,    0*2048+ 212,   17*2048+ 769,    0*2048+1117,
   0*2048+ 222,   13*2048+ 684,   19*2048+ 759,    0*2048+1118,
   0*2048+ 234,    6*2048+ 561,    1*2048+ 989,    0*2048+1119,
   0*2048+ 244,   17*2048+ 308,   32*2048+ 570,    0*2048+1120,
   0*2048+ 256,   29*2048+ 400,   14*2048+ 913,    0*2048+1121,
  28*2048+ 188,    0*2048+ 310,   22*2048+ 519,    0*2048+1123,
  42*2048+ 213,    0*2048+ 316,   32*2048+ 648,    0*2048+1124,
   0*2048+ 332,   35*2048+ 408,   27*2048+ 760,    0*2048+1125,
  40*2048+ 157,   36*2048+ 189,    0*2048+ 342,    0*2048+1126,
  43*2048+ 277,    0*2048+ 353,   21*2048+ 749,    0*2048+1127,
   0*2048+ 363,   28*2048+ 858,   43*2048+ 883,    0*2048+1128,
   0*2048+ 373,   41*2048+ 374,   11*2048+ 419,    0*2048+1129,
   0*2048+ 389,   10*2048+ 531,   23*2048+ 606,    0*2048+1130,
   0*2048+ 267,   15*2048+ 463,   31*2048+ 869,    0*2048+1131,
  14*2048+  91,    0*2048+ 278,   31*2048+ 562,    0*2048+1132,
  12*2048+ 103,   18*2048+ 134,    0*2048+ 288,    0*2048+1133,
  39*2048+  60,    0*2048+ 299,    1*2048+ 660,    0*2048+1134,
  19*2048+ 190,    0*2048+ 311,    6*2048+ 948,    0*2048+1135,
  36*2048+ 168,    0*2048+ 317,   18*2048+ 770,    0*2048+1136,
  38*2048+  92,    0*2048+ 333,   13*2048+ 364,    0*2048+1137,
   0*2048+ 343,   38*2048+ 771,    5*2048+ 949,    0*2048+1138,
   0*2048+ 354,   20*2048+ 540,   10*2048+ 870,    0*2048+1139,
   0*2048+ 365,   20*2048+ 571,    4*2048+ 572,    0*2048+1140,
   0*2048+ 375,   23*2048+ 596,   10*2048+ 649,    0*2048+1141,
  20*2048+ 124,    0*2048+ 390,   43*2048+ 409,    0*2048+1142,
  26*2048+  93,    0*2048+ 268,   32*2048+ 344,    0*2048+1143,
   0*2048+ 279,   11*2048+ 618,   31*2048+ 761,    0*2048+1144,
   0*2048+ 289,   14*2048+ 650,    7*2048+ 713,    0*2048+1145,
   0*2048+ 300,   10*2048+ 671,   40*2048+ 958,    0*2048+1146,
  35*2048+ 280,    0*2048+ 312,   24*2048+ 473,    0*2048+1147,
   0*2048+ 318,   10*2048+ 551,   11*2048+ 859,    0*2048+1148,
   0*2048+ 334,   26*2048+ 661,    1*2048+ 772,    0*2048+1149,
  25*2048+ 319,    0*2048+ 345,   17*2048+ 901,    0*2048+1150,
   0*2048+ 355,   13*2048+ 817,   19*2048+ 892,    0*2048+1151,
   2*2048+  68,    0*2048+ 366,    6*2048+ 694,    0*2048+1152,
   0*2048+ 376,   17*2048+ 441,   32*2048+ 702,    0*2048+1153,
   0*2048+ 391,   29*2048+ 532,   14*2048+1045,    0*2048+1154,
  28*2048+ 320,    0*2048+ 443,   22*2048+ 651,    0*2048+1156,
  42*2048+ 346,    0*2048+ 450,   32*2048+ 781,    0*2048+1157,
   0*2048+ 464,   35*2048+ 541,   27*2048+ 893,    0*2048+1158,
  40*2048+ 290,   36*2048+ 321,    0*2048+ 474,    0*2048+1159,
  43*2048+ 410,    0*2048+ 486,   21*2048+ 884,    0*2048+1160,
   0*2048+ 497,   28*2048+ 990,   43*2048+1015,    0*2048+1161,
   0*2048+ 508,   41*2048+ 509,   11*2048+ 552,    0*2048+1162,
   0*2048+ 521,   10*2048+ 663,   23*2048+ 738,    0*2048+1163,
   0*2048+ 401,   15*2048+ 597,   31*2048+1002,    0*2048+1164,
  14*2048+ 223,    0*2048+ 411,   31*2048+ 695,    0*2048+1165,
  12*2048+ 235,   18*2048+ 269,    0*2048+ 420,    0*2048+1166,
  39*2048+ 192,    0*2048+ 432,    1*2048+ 792,    0*2048+1167,
   7*2048+  26,   19*2048+ 322,    0*2048+ 444,    0*2048+1168,
  36*2048+ 301,    0*2048+ 451,   18*2048+ 902,    0*2048+1169,
  38*2048+ 224,    0*2048+ 465,   13*2048+ 498,    0*2048+1170,
   6*2048+  27,    0*2048+ 475,   38*2048+ 903,    0*2048+1171,
   0*2048+ 487,   20*2048+ 672,   10*2048+1003,    0*2048+1172,
   0*2048+ 499,   20*2048+ 703,    4*2048+ 704,    0*2048+1173,
   0*2048+ 510,   23*2048+ 728,   10*2048+ 782,    0*2048+1174,
  20*2048+ 257,    0*2048+ 522,   43*2048+ 542,    0*2048+1175,
  26*2048+ 225,    0*2048+ 402,   32*2048+ 476,    0*2048+1176,
   0*2048+ 412,   11*2048+ 750,   31*2048+ 894,    0*2048+1177,
   0*2048+ 421,   14*2048+ 783,    7*2048+ 847,    0*2048+1178,
  41*2048+  37,    0*2048+ 433,   10*2048+ 804,    0*2048+1179,
  35*2048+ 413,    0*2048+ 445,   24*2048+ 607,    0*2048+1180,
   0*2048+ 452,   10*2048+ 685,   11*2048+ 991,    0*2048+1181,
   0*2048+ 466,   26*2048+ 793,    1*2048+ 904,    0*2048+1182,
  25*2048+ 453,    0*2048+ 477,   17*2048+1034,    0*2048+1183,
   0*2048+ 488,   13*2048+ 950,   19*2048+1024,    0*2048+1184,
   2*2048+ 201,    0*2048+ 500,    6*2048+ 826,    0*2048+1185,
   0*2048+ 511,   17*2048+ 573,   32*2048+ 834,    0*2048+1186,
  15*2048+ 125,    0*2048+ 523,   29*2048+ 664,    0*2048+1187,
  28*2048+ 454,    0*2048+ 575,   22*2048+ 784,    0*2048+1189,
  42*2048+ 478,    0*2048+ 582,   32*2048+ 914,    0*2048+1190,
   0*2048+ 598,   35*2048+ 673,   27*2048+1025,    0*2048+1191,
  40*2048+ 422,   36*2048+ 455,    0*2048+ 608,    0*2048+1192,
  43*2048+ 543,    0*2048+ 619,   21*2048+1016,    0*2048+1193,
  29*2048+  69,   44*2048+  94,    0*2048+ 630,    0*2048+1194,
   0*2048+ 641,   41*2048+ 642,   11*2048+ 686,    0*2048+1195,
   0*2048+ 653,   10*2048+ 795,   23*2048+ 871,    0*2048+1196,
  32*2048+  82,    0*2048+ 533,   15*2048+ 729,    0*2048+1197,
  14*2048+ 356,    0*2048+ 544,   31*2048+ 827,    0*2048+1198,
  12*2048+ 367,   18*2048+ 403,    0*2048+ 553,    0*2048+1199,
  39*2048+ 324,    0*2048+ 564,    1*2048+ 925,    0*2048+1200,
   7*2048+ 159,   19*2048+ 456,    0*2048+ 576,    0*2048+1201,
  36*2048+ 434,    0*2048+ 583,   18*2048+1035,    0*2048+1202,
  38*2048+ 357,    0*2048+ 599,   13*2048+ 631,    0*2048+1203,
   6*2048+ 160,    0*2048+ 609,   38*2048+1036,    0*2048+1204,
  11*2048+  83,    0*2048+ 620,   20*2048+ 805,    0*2048+1205,
   0*2048+ 632,   20*2048+ 835,    4*2048+ 836,    0*2048+1206,
   0*2048+ 643,   23*2048+ 861,   10*2048+ 915,    0*2048+1207,
  20*2048+ 392,    0*2048+ 654,   43*2048+ 674,    0*2048+1208,
  26*2048+ 358,    0*2048+ 534,   32*2048+ 610,    0*2048+1209,
   0*2048+ 545,   11*2048+ 885,   31*2048+1026,    0*2048+1210,
   0*2048+ 554,   14*2048+ 916,    7*2048+ 982,    0*2048+1211,
  41*2048+ 169,    0*2048+ 565,   10*2048+ 936,    0*2048+1212,
  35*2048+ 546,    0*2048+ 577,   24*2048+ 739,    0*2048+1213,
  12*2048+  70,    0*2048+ 584,   10*2048+ 818,    0*2048+1214,
   0*2048+ 600,   26*2048+ 926,    1*2048+1037,    0*2048+1215,
  18*2048+ 114,   25*2048+ 585,    0*2048+ 611,    0*2048+1216,
  14*2048+  28,   20*2048+ 104,    0*2048+ 621,    0*2048+1217,
   2*2048+ 335,    0*2048+ 633,    6*2048+ 959,    0*2048+1218,
   0*2048+ 644,   17*2048+ 705,   32*2048+ 966,    0*2048+1219,
  15*2048+ 258,    0*2048+ 655,   29*2048+ 796,    0*2048+1220,
  28*2048+ 586,    0*2048+ 707,   22*2048+ 917,    0*2048+1222,
  42*2048+ 612,    0*2048+ 714,   32*2048+1046,    0*2048+1223,
  28*2048+ 105,    0*2048+ 730,   35*2048+ 806,    0*2048+1224,
  40*2048+ 555,   36*2048+ 587,    0*2048+ 740,    0*2048+1225,
  22*2048+  95,   43*2048+ 675,    0*2048+ 751,    0*2048+1226,
  29*2048+ 202,   44*2048+ 226,    0*2048+ 762,    0*2048+1227,
   0*2048+ 773,   41*2048+ 774,   11*2048+ 819,    0*2048+1228,
   0*2048+ 786,   10*2048+ 928,   23*2048+1004,    0*2048+1229,
  32*2048+ 215,    0*2048+ 665,   15*2048+ 862,    0*2048+1230,
  14*2048+ 489,    0*2048+ 676,   31*2048+ 960,    0*2048+1231,
  12*2048+ 501,   18*2048+ 535,    0*2048+ 687,    0*2048+1232,
   2*2048+   3,   39*2048+ 458,    0*2048+ 697,    0*2048+1233,
   7*2048+ 292,   19*2048+ 588,    0*2048+ 708,    0*2048+1234,
  19*2048+ 115,   36*2048+ 566,    0*2048+ 715,    0*2048+1235,
  38*2048+ 490,    0*2048+ 731,   13*2048+ 763,    0*2048+1236,
  39*2048+ 116,    6*2048+ 293,    0*2048+ 741,    0*2048+1237,
  11*2048+ 216,    0*2048+ 752,   20*2048+ 937,    0*2048+1238,
   0*2048+ 764,   20*2048+ 967,    4*2048+ 968,    0*2048+1239,
   0*2048+ 775,   23*2048+ 993,   10*2048+1047,    0*2048+1240,
  20*2048+ 524,    0*2048+ 787,   43*2048+ 807,    0*2048+1241,
  26*2048+ 491,    0*2048+ 666,   32*2048+ 742,    0*2048+1242,
  32*2048+ 106,    0*2048+ 677,   11*2048+1017,    0*2048+1243,
   8*2048+  62,    0*2048+ 688,   14*2048+1048,    0*2048+1244,
  11*2048+  16,   41*2048+ 302,    0*2048+ 698,    0*2048+1245,
  35*2048+ 678,    0*2048+ 709,   24*2048+ 872,    0*2048+1246,
  12*2048+ 203,    0*2048+ 716,   10*2048+ 951,    0*2048+1247,
  27*2048+   4,    2*2048+ 117,    0*2048+ 732,    0*2048+1248,
  18*2048+ 246,   25*2048+ 717,    0*2048+ 743,    0*2048+1249,
  14*2048+ 161,   20*2048+ 236,    0*2048+ 753,    0*2048+1250,
   7*2048+  38,    2*2048+ 467,    0*2048+ 765,    0*2048+1251,
  33*2048+  46,    0*2048+ 776,   17*2048+ 837,    0*2048+1252,
  15*2048+ 393,    0*2048+ 788,   29*2048+ 929,    0*2048+1253,
  28*2048+ 718,    0*2048+ 839,   22*2048+1049,    0*2048+1255,
  33*2048+ 126,   42*2048+ 744,    0*2048+ 848,    0*2048+1256,
  28*2048+ 237,    0*2048+ 863,   35*2048+ 938,    0*2048+1257,
  40*2048+ 689,   36*2048+ 719,    0*2048+ 873,    0*2048+1258,
  22*2048+ 227,   43*2048+ 808,    0*2048+ 886,    0*2048+1259,
  29*2048+ 336,   44*2048+ 359,    0*2048+ 895,    0*2048+1260,
   0*2048+ 905,   41*2048+ 906,   11*2048+ 952,    0*2048+1261,
  11*2048+   6,   24*2048+  84,    0*2048+ 919,    0*2048+1262,
  32*2048+ 348,    0*2048+ 797,   15*2048+ 994,    0*2048+1263,
  32*2048+  39,   14*2048+ 622,    0*2048+ 809,    0*2048+1264,
  12*2048+ 634,   18*2048+ 667,    0*2048+ 820,    0*2048+1265,
   2*2048+ 135,   39*2048+ 590,    0*2048+ 829,    0*2048+1266,
   7*2048+ 424,   19*2048+ 720,    0*2048+ 840,    0*2048+1267,
  19*2048+ 247,   36*2048+ 699,    0*2048+ 849,    0*2048+1268,
  38*2048+ 623,    0*2048+ 864,   13*2048+ 896,    0*2048+1269,
  39*2048+ 248,    6*2048+ 425,    0*2048+ 874,    0*2048+1270,
  21*2048+  17,   11*2048+ 349,    0*2048+ 887,    0*2048+1271,
  21*2048+  47,    5*2048+  48,    0*2048+ 897,    0*2048+1272,
  24*2048+  72,   11*2048+ 127,    0*2048+ 907,    0*2048+1273,
  20*2048+ 656,    0*2048+ 920,   43*2048+ 939,    0*2048+1274,
  26*2048+ 624,    0*2048+ 798,   32*2048+ 875,    0*2048+1275,
  12*2048+  96,   32*2048+ 238,    0*2048+ 810,    0*2048+1276,
  15*2048+ 128,    8*2048+ 194,    0*2048+ 821,    0*2048+1277,
  11*2048+ 150,   41*2048+ 435,    0*2048+ 830,    0*2048+1278,
  35*2048+ 811,    0*2048+ 841,   24*2048+1005,    0*2048+1279,
  11*2048+  29,   12*2048+ 337,    0*2048+ 850,    0*2048+1280,
  27*2048+ 136,    2*2048+ 249,    0*2048+ 865,    0*2048+1281,
  18*2048+ 378,   25*2048+ 851,    0*2048+ 876,    0*2048+1282,
  14*2048+ 294,   20*2048+ 368,    0*2048+ 888,    0*2048+1283,
   7*2048+ 170,    2*2048+ 601,    0*2048+ 898,    0*2048+1284,
  33*2048+ 179,    0*2048+ 908,   17*2048+ 969,    0*2048+1285,
  30*2048+   7,   15*2048+ 525,    0*2048+ 921,    0*2048+1286,
  23*2048+ 129,   28*2048+ 852,    0*2048+ 971,    0*2048+1288,
  33*2048+ 259,   42*2048+ 877,    0*2048+ 983,    0*2048+1289,
  36*2048+  18,   28*2048+ 369,    0*2048+ 995,    0*2048+1290,
  40*2048+ 822,   36*2048+ 853,    0*2048+1006,    0*2048+1291,
  22*2048+ 360,   43*2048+ 940,    0*2048+1018,    0*2048+1292,
  29*2048+ 468,   44*2048+ 492,    0*2048+1027,    0*2048+1293,
  12*2048+  30,    0*2048+1038,   41*2048+1039,    0*2048+1294,
  11*2048+ 138,   24*2048+ 217,    0*2048+1051,    0*2048+1295,
  16*2048+  73,   32*2048+ 480,    0*2048+ 930,    0*2048+1296,
  32*2048+ 171,   14*2048+ 754,    0*2048+ 941,    0*2048+1297,
  12*2048+ 766,   18*2048+ 799,    0*2048+ 953,    0*2048+1298,
   2*2048+ 270,   39*2048+ 722,    0*2048+ 962,    0*2048+1299,
   7*2048+ 557,   19*2048+ 854,    0*2048+ 972,    0*2048+1300,
  19*2048+ 379,   36*2048+ 831,    0*2048+ 984,    0*2048+1301,
  38*2048+ 755,    0*2048+ 996,   13*2048+1028,    0*2048+1302,
  39*2048+ 380,    6*2048+ 558,    0*2048+1007,    0*2048+1303,
  21*2048+ 151,   11*2048+ 481,    0*2048+1019,    0*2048+1304,
  21*2048+ 180,    5*2048+ 181,    0*2048+1029,    0*2048+1305,
  24*2048+ 205,   11*2048+ 260,    0*2048+1040,    0*2048+1306,
  44*2048+  19,   20*2048+ 789,    0*2048+1052,    0*2048+1307,
  26*2048+ 756,    0*2048+ 931,   32*2048+1008,    0*2048+1308,
  12*2048+ 228,   32*2048+ 370,    0*2048+ 942,    0*2048+1309,
  15*2048+ 261,    8*2048+ 326,    0*2048+ 954,    0*2048+1310,
  11*2048+ 283,   41*2048+ 567,    0*2048+ 963,    0*2048+1311,
  25*2048+  85,   35*2048+ 943,    0*2048+ 973,    0*2048+1312,
  11*2048+ 162,   12*2048+ 469,    0*2048+ 985,    0*2048+1313,
  27*2048+ 271,    2*2048+ 381,    0*2048+ 997,    0*2048+1314,
  18*2048+ 513,   25*2048+ 986,    0*2048+1009,    0*2048+1315,
  14*2048+ 426,   20*2048+ 502,    0*2048+1020,    0*2048+1316,
   7*2048+ 303,    2*2048+ 733,    0*2048+1030,    0*2048+1317,
  18*2048+  49,   33*2048+ 313,    0*2048+1041,    0*2048+1318,
  30*2048+ 139,   15*2048+ 657,    0*2048+1053,    0*2048+1319,
   0*2048+  33,   20*2048+  42,    7*2048+ 120,   27*2048+ 264,   33*2048+ 329,   15*2048+ 448,   10*2048+ 538,   18*2048+ 802,    5*2048+ 814,   35*2048+ 844,   43*2048+ 868,    4*2048+1033,    0*2048+1056,
   5*2048+ 113,    0*2048+ 165,   20*2048+ 175,    7*2048+ 253,   27*2048+ 398,   33*2048+ 461,   15*2048+ 580,   10*2048+ 670,   18*2048+ 934,    5*2048+ 947,   35*2048+ 979,   43*2048+1001,    0*2048+1089,
  19*2048+  14,    6*2048+  25,   36*2048+  59,   44*2048+  81,    5*2048+ 245,    0*2048+ 298,   20*2048+ 309,    7*2048+ 388,   27*2048+ 530,   33*2048+ 595,   15*2048+ 712,   10*2048+ 803,    0*2048+1122,
  19*2048+ 148,    6*2048+ 158,   36*2048+ 191,   44*2048+ 214,    5*2048+ 377,    0*2048+ 431,   20*2048+ 442,    7*2048+ 520,   27*2048+ 662,   33*2048+ 727,   15*2048+ 846,   10*2048+ 935,    0*2048+1155,
  11*2048+  15,   19*2048+ 281,    6*2048+ 291,   36*2048+ 323,   44*2048+ 347,    5*2048+ 512,    0*2048+ 563,   20*2048+ 574,    7*2048+ 652,   27*2048+ 794,   33*2048+ 860,   15*2048+ 981,    0*2048+1188,
  16*2048+  61,   11*2048+ 149,   19*2048+ 414,    6*2048+ 423,   36*2048+ 457,   44*2048+ 479,    5*2048+ 645,    0*2048+ 696,   20*2048+ 706,    7*2048+ 785,   27*2048+ 927,   33*2048+ 992,    0*2048+1221,
  28*2048+   5,   34*2048+  71,   16*2048+ 193,   11*2048+ 282,   19*2048+ 547,    6*2048+ 556,   36*2048+ 589,   44*2048+ 613,    5*2048+ 777,    0*2048+ 828,   20*2048+ 838,    7*2048+ 918,    0*2048+1254,
  28*2048+ 137,   34*2048+ 204,   16*2048+ 325,   11*2048+ 415,   19*2048+ 679,    6*2048+ 690,   36*2048+ 721,   44*2048+ 745,    5*2048+ 909,    0*2048+ 961,   20*2048+ 970,    7*2048+1050,    0*2048+1287,

   0*2048+  10,    0*2048+  21,    0*2048+1280,
   0*2048+  22,    0*2048+  34,    0*2048+1281,
   0*2048+  35,    0*2048+  46,    0*2048+1282,
   0*2048+  47,    0*2048+  58,    0*2048+1283,
   0*2048+  59,    0*2048+  71,    0*2048+1284,
   0*2048+  72,    0*2048+  84,    0*2048+1285,
   0*2048+  85,    0*2048+  97,    0*2048+1286,
   0*2048+  98,    0*2048+ 110,    0*2048+1287,
   0*2048+ 111,    0*2048+ 123,    0*2048+1288,
   0*2048+ 124,    0*2048+ 135,    0*2048+1289,
   0*2048+ 136,    0*2048+ 146,    0*2048+1290,
   0*2048+ 147,    0*2048+ 159,    0*2048+1291,
   0*2048+ 160,    0*2048+ 171,    0*2048+1292,
   0*2048+ 172,    0*2048+ 183,    0*2048+1293,
   0*2048+ 184,    0*2048+ 196,    0*2048+1294,
   0*2048+ 197,    0*2048+ 209,    0*2048+1295,
   0*2048+ 210,    0*2048+ 222,    0*2048+1296,
   0*2048+ 223,    0*2048+ 235,    0*2048+1297,
   0*2048+ 236,    0*2048+ 248,    0*2048+1298,
   0*2048+ 249,    0*2048+ 260,    0*2048+1299,
   0*2048+ 261,    0*2048+ 271,    0*2048+1300,
   0*2048+ 272,    0*2048+ 284,    0*2048+1301,
   0*2048+ 285,    0*2048+ 296,    0*2048+1302,
   0*2048+ 297,    0*2048+ 308,    0*2048+1303,
   0*2048+ 309,    0*2048+ 321,    0*2048+1304,
   0*2048+ 322,    0*2048+ 334,    0*2048+1305,
   0*2048+ 335,    0*2048+ 347,    0*2048+1306,
   0*2048+ 348,    0*2048+ 360,    0*2048+1307,
   0*2048+ 361,    0*2048+ 373,    0*2048+1308,
   0*2048+ 374,    0*2048+ 385,    0*2048+1309,
   0*2048+ 386,    0*2048+ 396,    0*2048+1310,
   0*2048+ 397,    0*2048+ 409,    0*2048+1311,
   0*2048+ 410,    0*2048+ 421,    0*2048+1312,
   0*2048+ 422,    0*2048+ 433,    0*2048+1313,
   0*2048+ 434,    0*2048+ 446,    0*2048+1314,
   0*2048+ 447,    0*2048+ 459,    0*2048+1315,
   0*2048+ 460,    0*2048+ 472,    0*2048+1316,
   0*2048+ 473,    0*2048+ 485,    0*2048+1317,
   0*2048+ 486,    0*2048+ 498,    0*2048+1318,
   0*2048+ 499,    0*2048+ 510,    0*2048+1319,
   0*2048+ 511,    0*2048+ 521,    0*2048+1320,
   0*2048+ 522,    0*2048+ 534,    0*2048+1321,
   0*2048+ 535,    0*2048+ 546,    0*2048+1322,
   0*2048+ 547,    0*2048+ 558,    0*2048+1323,
   0*2048+ 559,    0*2048+ 571,    0*2048+1324,
   0*2048+ 572,    0*2048+ 584,    0*2048+1325,
   0*2048+ 585,    0*2048+ 597,    0*2048+1326,
   0*2048+ 598,    0*2048+ 610,    0*2048+1327,
   0*2048+ 611,    0*2048+ 623,    0*2048+1328,
   0*2048+ 624,    0*2048+ 635,    0*2048+1329,
   0*2048+ 636,    0*2048+ 646,    0*2048+1330,
   0*2048+ 647,    0*2048+ 659,    0*2048+1331,
   0*2048+ 660,    0*2048+ 671,    0*2048+1332,
   0*2048+ 672,    0*2048+ 683,    0*2048+1333,
   0*2048+ 684,    0*2048+ 696,    0*2048+1334,
   0*2048+ 697,    0*2048+ 709,    0*2048+1335,
   0*2048+ 710,    0*2048+ 722,    0*2048+1336,
   0*2048+ 723,    0*2048+ 735,    0*2048+1337,
   0*2048+ 736,    0*2048+ 748,    0*2048+1338,
   0*2048+ 749,    0*2048+ 760,    0*2048+1339,
   0*2048+ 761,    0*2048+ 771,    0*2048+1340,
   0*2048+ 772,    0*2048+ 784,    0*2048+1341,
   0*2048+ 785,    0*2048+ 796,    0*2048+1342,
   0*2048+ 797,    0*2048+ 808,    0*2048+1343,
   0*2048+ 809,    0*2048+ 821,    0*2048+1344,
   0*2048+ 822,    0*2048+ 834,    0*2048+1345,
   0*2048+ 835,    0*2048+ 847,    0*2048+1346,
   0*2048+ 848,    0*2048+ 860,    0*2048+1347,
   0*2048+ 861,    0*2048+ 873,    0*2048+1348,
   0*2048+ 874,    0*2048+ 885,    0*2048+1349,
   0*2048+ 886,    0*2048+ 896,    0*2048+1350,
   0*2048+ 897,    0*2048+ 909,    0*2048+1351,
   0*2048+ 910,    0*2048+ 921,    0*2048+1352,
   0*2048+ 922,    0*2048+ 933,    0*2048+1353,
   0*2048+ 934,    0*2048+ 946,    0*2048+1354,
   0*2048+ 947,    0*2048+ 959,    0*2048+1355,
   0*2048+ 960,    0*2048+ 972,    0*2048+1356,
   0*2048+ 973,    0*2048+ 985,    0*2048+1357,
   0*2048+ 986,    0*2048+ 998,    0*2048+1358,
   1*2048+  11,    0*2048+ 999,    0*2048+1359,
   0*2048+  60,   11*2048+ 198,   19*2048+ 560,    0*2048+1000,
   0*2048+  73,   31*2048+ 161,    2*2048+ 298,    0*2048+1001,
   0*2048+  86,   40*2048+ 125,    2*2048+ 648,    0*2048+1002,
   9*2048+  87,    0*2048+  99,   16*2048+ 737,    0*2048+1003,
   0*2048+ 112,    7*2048+ 649,   42*2048+ 849,    0*2048+1004,
   0*2048+   0,   33*2048+ 286,   24*2048+ 336,    0*2048+1005,
   0*2048+  12,   33*2048+ 685,    2*2048+ 875,    0*2048+1006,
   0*2048+  23,   25*2048+ 310,   34*2048+ 923,    0*2048+1007,
   0*2048+  36,    3*2048+ 536,   37*2048+ 987,    0*2048+1008,
   0*2048+  48,   36*2048+ 113,   10*2048+ 773,    0*2048+1009,
   0*2048+  61,   26*2048+ 375,    4*2048+ 698,    0*2048+1010,
   0*2048+  74,   25*2048+ 423,   28*2048+ 573,    0*2048+1011,
   0*2048+  88,   25*2048+ 850,   11*2048+ 887,    0*2048+1012,
   0*2048+ 100,   44*2048+ 273,   38*2048+ 851,    0*2048+1013,
   0*2048+ 114,   17*2048+ 762,    3*2048+ 836,    0*2048+1014,
   0*2048+   1,   28*2048+ 398,   14*2048+ 961,    0*2048+1015,
  41*2048+   2,    0*2048+  13,   22*2048+ 500,    0*2048+1016,
   0*2048+  24,    4*2048+ 137,   28*2048+ 852,    0*2048+1017,
   0*2048+  37,    5*2048+ 810,   31*2048+ 898,    0*2048+1018,
   0*2048+  49,   12*2048+ 974,   30*2048+ 988,    0*2048+1019,
   0*2048+  62,   17*2048+ 287,    4*2048+ 288,    0*2048+1020,
   0*2048+  75,    1*2048+ 173,    2*2048+ 948,    0*2048+1021,
   0*2048+  89,    1*2048+ 512,   32*2048+ 738,    0*2048+1022,
   0*2048+ 101,   34*2048+ 673,   18*2048+ 711,    0*2048+1023,
   0*2048+ 115,   23*2048+ 185,   26*2048+ 448,    0*2048+1024,
   0*2048+   3,    9*2048+  25,   19*2048+ 798,    0*2048+1025,
   0*2048+  14,   23*2048+ 513,   34*2048+ 586,    0*2048+1026,
   0*2048+  26,   20*2048+ 126,   33*2048+ 763,    0*2048+1027,
   0*2048+  38,   41*2048+  39,   21*2048+ 650,    0*2048+1028,
   0*2048+  50,    2*2048+ 102,   13*2048+ 739,    0*2048+1029,
   3*2048+  40,    0*2048+  63,   38*2048+ 424,    0*2048+1030,
   0*2048+  76,   43*2048+ 250,   11*2048+ 811,    0*2048+1031,
   0*2048+  90,   25*2048+ 612,   21*2048+ 823,    0*2048+1032,
   7*2048+  77,    0*2048+ 103,   17*2048+ 837,    0*2048+1033,
   0*2048+ 116,   44*2048+ 311,   14*2048+ 599,    0*2048+1034,
   0*2048+ 186,   11*2048+ 323,   19*2048+ 686,    0*2048+1035,
   0*2048+ 199,   31*2048+ 289,    2*2048+ 425,    0*2048+1036,
   0*2048+ 211,   40*2048+ 251,    2*2048+ 774,    0*2048+1037,
   9*2048+ 212,    0*2048+ 224,   16*2048+ 862,    0*2048+1038,
   0*2048+ 237,    7*2048+ 775,   42*2048+ 975,    0*2048+1039,
   0*2048+ 127,   33*2048+ 411,   24*2048+ 461,    0*2048+1040,
   3*2048+   4,    0*2048+ 138,   33*2048+ 812,    0*2048+1041,
  35*2048+  51,    0*2048+ 148,   25*2048+ 435,    0*2048+1042,
  38*2048+ 117,    0*2048+ 162,    3*2048+ 661,    0*2048+1043,
   0*2048+ 174,   36*2048+ 238,   10*2048+ 899,    0*2048+1044,
   0*2048+ 187,   26*2048+ 501,    4*2048+ 824,    0*2048+1045,
   0*2048+ 200,   25*2048+ 548,   28*2048+ 699,    0*2048+1046,
  12*2048+  15,    0*2048+ 213,   25*2048+ 976,    0*2048+1047,
   0*2048+ 225,   44*2048+ 399,   38*2048+ 977,    0*2048+1048,
   0*2048+ 239,   17*2048+ 888,    3*2048+ 962,    0*2048+1049,
  15*2048+  91,    0*2048+ 128,   28*2048+ 523,    0*2048+1050,
  41*2048+ 129,    0*2048+ 139,   22*2048+ 625,    0*2048+1051,
   0*2048+ 149,    4*2048+ 262,   28*2048+ 978,    0*2048+1052,
  32*2048+  27,    0*2048+ 163,    5*2048+ 935,    0*2048+1053,
  13*2048+ 104,   31*2048+ 118,    0*2048+ 175,    0*2048+1054,
   0*2048+ 188,   17*2048+ 412,    4*2048+ 413,    0*2048+1055,
   3*2048+  78,    0*2048+ 201,    1*2048+ 299,    0*2048+1056,
   0*2048+ 214,    1*2048+ 637,   32*2048+ 863,    0*2048+1057,
   0*2048+ 226,   34*2048+ 799,   18*2048+ 838,    0*2048+1058,
   0*2048+ 240,   23*2048+ 312,   26*2048+ 574,    0*2048+1059,
   0*2048+ 130,    9*2048+ 150,   19*2048+ 924,    0*2048+1060,
   0*2048+ 140,   23*2048+ 638,   34*2048+ 712,    0*2048+1061,
   0*2048+ 151,   20*2048+ 252,   33*2048+ 889,    0*2048+1062,
   0*2048+ 164,   41*2048+ 165,   21*2048+ 776,    0*2048+1063,
   0*2048+ 176,    2*2048+ 227,   13*2048+ 864,    0*2048+1064,
   3*2048+ 166,    0*2048+ 189,   38*2048+ 549,    0*2048+1065,
   0*2048+ 202,   43*2048+ 376,   11*2048+ 936,    0*2048+1066,
   0*2048+ 215,   25*2048+ 740,   21*2048+ 949,    0*2048+1067,
   7*2048+ 203,    0*2048+ 228,   17*2048+ 963,    0*2048+1068,
   0*2048+ 241,   44*2048+ 436,   14*2048+ 724,    0*2048+1069,
   0*2048+ 313,   11*2048+ 449,   19*2048+ 813,    0*2048+1070,
   0*2048+ 324,   31*2048+ 414,    2*2048+ 550,    0*2048+1071,
   0*2048+ 337,   40*2048+ 377,    2*2048+ 900,    0*2048+1072,
   9*2048+ 338,    0*2048+ 349,   16*2048+ 989,    0*2048+1073,
  43*2048+ 105,    0*2048+ 362,    7*2048+ 901,    0*2048+1074,
   0*2048+ 253,   33*2048+ 537,   24*2048+ 587,    0*2048+1075,
   3*2048+ 131,    0*2048+ 263,   33*2048+ 937,    0*2048+1076,
  35*2048+ 177,    0*2048+ 274,   25*2048+ 561,    0*2048+1077,
  38*2048+ 242,    0*2048+ 290,    3*2048+ 786,    0*2048+1078,
  11*2048+  28,    0*2048+ 300,   36*2048+ 363,    0*2048+1079,
   0*2048+ 314,   26*2048+ 626,    4*2048+ 950,    0*2048+1080,
   0*2048+ 325,   25*2048+ 674,   28*2048+ 825,    0*2048+1081,
  26*2048+ 106,   12*2048+ 141,    0*2048+ 339,    0*2048+1082,
  39*2048+ 107,    0*2048+ 350,   44*2048+ 524,    0*2048+1083,
  18*2048+  16,    4*2048+  92,    0*2048+ 364,    0*2048+1084,
  15*2048+ 216,    0*2048+ 254,   28*2048+ 651,    0*2048+1085,
  41*2048+ 255,    0*2048+ 264,   22*2048+ 750,    0*2048+1086,
  29*2048+ 108,    0*2048+ 275,    4*2048+ 387,    0*2048+1087,
   6*2048+  64,   32*2048+ 152,    0*2048+ 291,    0*2048+1088,
  13*2048+ 229,   31*2048+ 243,    0*2048+ 301,    0*2048+1089,
   0*2048+ 315,   17*2048+ 538,    4*2048+ 539,    0*2048+1090,
   3*2048+ 204,    0*2048+ 326,    1*2048+ 426,    0*2048+1091,
   0*2048+ 340,    1*2048+ 764,   32*2048+ 990,    0*2048+1092,
   0*2048+ 351,   34*2048+ 925,   18*2048+ 964,    0*2048+1093,
   0*2048+ 365,   23*2048+ 437,   26*2048+ 700,    0*2048+1094,
  20*2048+  52,    0*2048+ 256,    9*2048+ 276,    0*2048+1095,
   0*2048+ 265,   23*2048+ 765,   34*2048+ 839,    0*2048+1096,
  34*2048+  17,    0*2048+ 277,   20*2048+ 378,    0*2048+1097,
   0*2048+ 292,   41*2048+ 293,   21*2048+ 902,    0*2048+1098,
   0*2048+ 302,    2*2048+ 352,   13*2048+ 991,    0*2048+1099,
   3*2048+ 294,    0*2048+ 316,   38*2048+ 675,    0*2048+1100,
  12*2048+  65,    0*2048+ 327,   43*2048+ 502,    0*2048+1101,
  22*2048+  79,    0*2048+ 341,   25*2048+ 865,    0*2048+1102,
  18*2048+  93,    7*2048+ 328,    0*2048+ 353,    0*2048+1103,
   0*2048+ 366,   44*2048+ 562,   14*2048+ 853,    0*2048+1104,
   0*2048+ 438,   11*2048+ 575,   19*2048+ 938,    0*2048+1105,
   0*2048+ 450,   31*2048+ 540,    2*2048+ 676,    0*2048+1106,
   3*2048+  29,    0*2048+ 462,   40*2048+ 503,    0*2048+1107,
  17*2048+ 119,    9*2048+ 463,    0*2048+ 474,    0*2048+1108,
   8*2048+  30,   43*2048+ 230,    0*2048+ 487,    0*2048+1109,
   0*2048+ 379,   33*2048+ 662,   24*2048+ 713,    0*2048+1110,
  34*2048+  66,    3*2048+ 257,    0*2048+ 388,    0*2048+1111,
  35*2048+ 303,    0*2048+ 400,   25*2048+ 687,    0*2048+1112,
  38*2048+ 367,    0*2048+ 415,    3*2048+ 911,    0*2048+1113,
  11*2048+ 153,    0*2048+ 427,   36*2048+ 488,    0*2048+1114,
   5*2048+  80,    0*2048+ 439,   26*2048+ 751,    0*2048+1115,
   0*2048+ 451,   25*2048+ 800,   28*2048+ 951,    0*2048+1116,
  26*2048+ 231,   12*2048+ 266,    0*2048+ 464,    0*2048+1117,
  39*2048+ 232,    0*2048+ 475,   44*2048+ 652,    0*2048+1118,
  18*2048+ 142,    4*2048+ 217,    0*2048+ 489,    0*2048+1119,
  15*2048+ 342,    0*2048+ 380,   28*2048+ 777,    0*2048+1120,
  41*2048+ 381,    0*2048+ 389,   22*2048+ 876,    0*2048+1121,
  29*2048+ 233,    0*2048+ 401,    4*2048+ 514,    0*2048+1122,
   6*2048+ 190,   32*2048+ 278,    0*2048+ 416,    0*2048+1123,
  13*2048+ 354,   31*2048+ 368,    0*2048+ 428,    0*2048+1124,
   0*2048+ 440,   17*2048+ 663,    4*2048+ 664,    0*2048+1125,
   3*2048+ 329,    0*2048+ 452,    1*2048+ 551,    0*2048+1126,
  33*2048+ 120,    0*2048+ 465,    1*2048+ 890,    0*2048+1127,
  35*2048+  53,   19*2048+  94,    0*2048+ 476,    0*2048+1128,
   0*2048+ 490,   23*2048+ 563,   26*2048+ 826,    0*2048+1129,
  20*2048+ 178,    0*2048+ 382,    9*2048+ 402,    0*2048+1130,
   0*2048+ 390,   23*2048+ 891,   34*2048+ 965,    0*2048+1131,
  34*2048+ 143,    0*2048+ 403,   20*2048+ 504,    0*2048+1132,
  22*2048+  31,    0*2048+ 417,   41*2048+ 418,    0*2048+1133,
  14*2048+ 121,    0*2048+ 429,    2*2048+ 477,    0*2048+1134,
   3*2048+ 419,    0*2048+ 441,   38*2048+ 801,    0*2048+1135,
  12*2048+ 191,    0*2048+ 453,   43*2048+ 627,    0*2048+1136,
  22*2048+ 205,    0*2048+ 466,   25*2048+ 992,    0*2048+1137,
  18*2048+ 218,    7*2048+ 454,    0*2048+ 478,    0*2048+1138,
   0*2048+ 491,   44*2048+ 688,   14*2048+ 979,    0*2048+1139,
  20*2048+  67,    0*2048+ 564,   11*2048+ 701,    0*2048+1140,
   0*2048+ 576,   31*2048+ 665,    2*2048+ 802,    0*2048+1141,
   3*2048+ 154,    0*2048+ 588,   40*2048+ 628,    0*2048+1142,
  17*2048+ 244,    9*2048+ 589,    0*2048+ 600,    0*2048+1143,
   8*2048+ 155,   43*2048+ 355,    0*2048+ 613,    0*2048+1144,
   0*2048+ 505,   33*2048+ 787,   24*2048+ 840,    0*2048+1145,
  34*2048+ 192,    3*2048+ 383,    0*2048+ 515,    0*2048+1146,
  35*2048+ 430,    0*2048+ 525,   25*2048+ 814,    0*2048+1147,
   4*2048+  41,   38*2048+ 492,    0*2048+ 541,    0*2048+1148,
  11*2048+ 279,    0*2048+ 552,   36*2048+ 614,    0*2048+1149,
   5*2048+ 206,    0*2048+ 565,   26*2048+ 877,    0*2048+1150,
  29*2048+  81,    0*2048+ 577,   25*2048+ 926,    0*2048+1151,
  26*2048+ 356,   12*2048+ 391,    0*2048+ 590,    0*2048+1152,
  39*2048+ 357,    0*2048+ 601,   44*2048+ 778,    0*2048+1153,
  18*2048+ 267,    4*2048+ 343,    0*2048+ 615,    0*2048+1154,
  15*2048+ 467,    0*2048+ 506,   28*2048+ 903,    0*2048+1155,
  23*2048+   5,   41*2048+ 507,    0*2048+ 516,    0*2048+1156,
  29*2048+ 358,    0*2048+ 526,    4*2048+ 639,    0*2048+1157,
   6*2048+ 317,   32*2048+ 404,    0*2048+ 542,    0*2048+1158,
  13*2048+ 479,   31*2048+ 493,    0*2048+ 553,    0*2048+1159,
   0*2048+ 566,   17*2048+ 788,    4*2048+ 789,    0*2048+1160,
   3*2048+ 455,    0*2048+ 578,    1*2048+ 677,    0*2048+1161,
   2*2048+  18,   33*2048+ 245,    0*2048+ 591,    0*2048+1162,
  35*2048+ 179,   19*2048+ 219,    0*2048+ 602,    0*2048+1163,
   0*2048+ 616,   23*2048+ 689,   26*2048+ 952,    0*2048+1164,
  20*2048+ 304,    0*2048+ 508,    9*2048+ 527,    0*2048+1165,
  24*2048+  19,   35*2048+  95,    0*2048+ 517,    0*2048+1166,
  34*2048+ 268,    0*2048+ 528,   20*2048+ 629,    0*2048+1167,
  22*2048+ 156,    0*2048+ 543,   41*2048+ 544,    0*2048+1168,
  14*2048+ 246,    0*2048+ 554,    2*2048+ 603,    0*2048+1169,
   3*2048+ 545,    0*2048+ 567,   38*2048+ 927,    0*2048+1170,
  12*2048+ 318,    0*2048+ 579,   43*2048+ 752,    0*2048+1171,
  26*2048+ 122,   22*2048+ 330,    0*2048+ 592,    0*2048+1172,
  18*2048+ 344,    7*2048+ 580,    0*2048+ 604,    0*2048+1173,
  15*2048+ 109,    0*2048+ 617,   44*2048+ 815,    0*2048+1174,
  20*2048+ 193,    0*2048+ 690,   11*2048+ 827,    0*2048+1175,
   0*2048+ 702,   31*2048+ 790,    2*2048+ 928,    0*2048+1176,
   3*2048+ 280,    0*2048+ 714,   40*2048+ 753,    0*2048+1177,
  17*2048+ 369,    9*2048+ 715,    0*2048+ 725,    0*2048+1178,
   8*2048+ 281,   43*2048+ 480,    0*2048+ 741,    0*2048+1179,
   0*2048+ 630,   33*2048+ 912,   24*2048+ 966,    0*2048+1180,
  34*2048+ 319,    3*2048+ 509,    0*2048+ 640,    0*2048+1181,
  35*2048+ 555,    0*2048+ 653,   25*2048+ 939,    0*2048+1182,
   4*2048+ 167,   38*2048+ 618,    0*2048+ 666,    0*2048+1183,
  11*2048+ 405,    0*2048+ 678,   36*2048+ 742,    0*2048+1184,
  27*2048+   6,    5*2048+ 331,    0*2048+ 691,    0*2048+1185,
  26*2048+  54,   29*2048+ 207,    0*2048+ 703,    0*2048+1186,
  26*2048+ 481,   12*2048+ 518,    0*2048+ 716,    0*2048+1187,
  39*2048+ 482,    0*2048+ 726,   44*2048+ 904,    0*2048+1188,
  18*2048+ 392,    4*2048+ 468,    0*2048+ 743,    0*2048+1189,
  29*2048+  32,   15*2048+ 593,    0*2048+ 631,    0*2048+1190,
  23*2048+ 132,   41*2048+ 632,    0*2048+ 641,    0*2048+1191,
  29*2048+ 483,    0*2048+ 654,    4*2048+ 766,    0*2048+1192,
   6*2048+ 442,   32*2048+ 529,    0*2048+ 667,    0*2048+1193,
  13*2048+ 605,   31*2048+ 619,    0*2048+ 679,    0*2048+1194,
   0*2048+ 692,   17*2048+ 913,    4*2048+ 914,    0*2048+1195,
   3*2048+ 581,    0*2048+ 704,    1*2048+ 803,    0*2048+1196,
   2*2048+ 144,   33*2048+ 370,    0*2048+ 717,    0*2048+1197,
  35*2048+ 305,   19*2048+ 345,    0*2048+ 727,    0*2048+1198,
  27*2048+  82,    0*2048+ 744,   23*2048+ 816,    0*2048+1199,
  20*2048+ 431,    0*2048+ 633,    9*2048+ 655,    0*2048+1200,
  24*2048+ 145,   35*2048+ 220,    0*2048+ 642,    0*2048+1201,
  34*2048+ 393,    0*2048+ 656,   20*2048+ 754,    0*2048+1202,
  22*2048+ 282,    0*2048+ 668,   41*2048+ 669,    0*2048+1203,
  14*2048+ 371,    0*2048+ 680,    2*2048+ 728,    0*2048+1204,
  39*2048+  55,    3*2048+ 670,    0*2048+ 693,    0*2048+1205,
  12*2048+ 443,    0*2048+ 705,   43*2048+ 878,    0*2048+1206,
  26*2048+ 247,   22*2048+ 456,    0*2048+ 718,    0*2048+1207,
  18*2048+ 469,    7*2048+ 706,    0*2048+ 729,    0*2048+1208,
  15*2048+ 234,    0*2048+ 745,   44*2048+ 940,    0*2048+1209,
  20*2048+ 320,    0*2048+ 817,   11*2048+ 953,    0*2048+1210,
   3*2048+  56,    0*2048+ 828,   31*2048+ 915,    0*2048+1211,
   3*2048+ 406,    0*2048+ 841,   40*2048+ 879,    0*2048+1212,
  17*2048+ 494,    9*2048+ 842,    0*2048+ 854,    0*2048+1213,
   8*2048+ 407,   43*2048+ 606,    0*2048+ 866,    0*2048+1214,
  34*2048+  42,   25*2048+  96,    0*2048+ 755,    0*2048+1215,
  34*2048+ 444,    3*2048+ 634,    0*2048+ 767,    0*2048+1216,
  26*2048+  68,   35*2048+ 681,    0*2048+ 779,    0*2048+1217,
   4*2048+ 295,   38*2048+ 746,    0*2048+ 791,    0*2048+1218,
  11*2048+ 530,    0*2048+ 804,   36*2048+ 867,    0*2048+1219,
  27*2048+ 133,    5*2048+ 457,    0*2048+ 818,    0*2048+1220,
  26*2048+ 180,   29*2048+ 332,    0*2048+ 829,    0*2048+1221,
  26*2048+ 607,   12*2048+ 643,    0*2048+ 843,    0*2048+1222,
  45*2048+  33,   39*2048+ 608,    0*2048+ 855,    0*2048+1223,
  18*2048+ 519,    4*2048+ 594,    0*2048+ 868,    0*2048+1224,
  29*2048+ 157,   15*2048+ 719,    0*2048+ 756,    0*2048+1225,
  23*2048+ 258,   41*2048+ 757,    0*2048+ 768,    0*2048+1226,
  29*2048+ 609,    0*2048+ 780,    4*2048+ 892,    0*2048+1227,
   6*2048+ 568,   32*2048+ 657,    0*2048+ 792,    0*2048+1228,
  13*2048+ 730,   31*2048+ 747,    0*2048+ 805,    0*2048+1229,
  18*2048+  43,    5*2048+  44,    0*2048+ 819,    0*2048+1230,
   3*2048+ 707,    0*2048+ 830,    1*2048+ 929,    0*2048+1231,
   2*2048+ 269,   33*2048+ 495,    0*2048+ 844,    0*2048+1232,
  35*2048+ 432,   19*2048+ 470,    0*2048+ 856,    0*2048+1233,
  27*2048+ 208,    0*2048+ 869,   23*2048+ 941,    0*2048+1234,
  20*2048+ 556,    0*2048+ 758,    9*2048+ 781,    0*2048+1235,
  24*2048+ 270,   35*2048+ 346,    0*2048+ 769,    0*2048+1236,
  34*2048+ 520,    0*2048+ 782,   20*2048+ 880,    0*2048+1237,
  22*2048+ 408,    0*2048+ 793,   41*2048+ 794,    0*2048+1238,
  14*2048+ 496,    0*2048+ 806,    2*2048+ 857,    0*2048+1239,
  39*2048+ 181,    3*2048+ 795,    0*2048+ 820,    0*2048+1240,
  44*2048+   7,   12*2048+ 569,    0*2048+ 831,    0*2048+1241,
  26*2048+ 372,   22*2048+ 582,    0*2048+ 845,    0*2048+1242,
  18*2048+ 595,    7*2048+ 832,    0*2048+ 858,    0*2048+1243,
  45*2048+  69,   15*2048+ 359,    0*2048+ 870,    0*2048+1244,
  12*2048+  83,   20*2048+ 445,    0*2048+ 942,    0*2048+1245,
  32*2048+  45,    3*2048+ 182,    0*2048+ 954,    0*2048+1246,
  41*2048+   8,    3*2048+ 531,    0*2048+ 967,    0*2048+1247,
  17*2048+ 620,    9*2048+ 968,    0*2048+ 980,    0*2048+1248,
   8*2048+ 532,   43*2048+ 731,    0*2048+ 993,    0*2048+1249,
  34*2048+ 168,   25*2048+ 221,    0*2048+ 881,    0*2048+1250,
  34*2048+ 570,    3*2048+ 759,    0*2048+ 893,    0*2048+1251,
  26*2048+ 194,   35*2048+ 807,    0*2048+ 905,    0*2048+1252,
   4*2048+ 420,   38*2048+ 871,    0*2048+ 916,    0*2048+1253,
  11*2048+ 658,    0*2048+ 930,   36*2048+ 994,    0*2048+1254,
  27*2048+ 259,    5*2048+ 583,    0*2048+ 943,    0*2048+1255,
  26*2048+ 306,   29*2048+ 458,    0*2048+ 955,    0*2048+1256,
  26*2048+ 732,   12*2048+ 770,    0*2048+ 969,    0*2048+1257,
  45*2048+ 158,   39*2048+ 733,    0*2048+ 981,    0*2048+1258,
  18*2048+ 644,    4*2048+ 720,    0*2048+ 995,    0*2048+1259,
  29*2048+ 283,   15*2048+ 846,    0*2048+ 882,    0*2048+1260,
  23*2048+ 384,   41*2048+ 883,    0*2048+ 894,    0*2048+1261,
   5*2048+  20,   29*2048+ 734,    0*2048+ 906,    0*2048+1262,
   6*2048+ 694,   32*2048+ 783,    0*2048+ 917,    0*2048+1263,
  13*2048+ 859,   31*2048+ 872,    0*2048+ 931,    0*2048+1264,
  18*2048+ 169,    5*2048+ 170,    0*2048+ 944,    0*2048+1265,
   2*2048+  57,    3*2048+ 833,    0*2048+ 956,    0*2048+1266,
   2*2048+ 394,   33*2048+ 621,    0*2048+ 970,    0*2048+1267,
  35*2048+ 557,   19*2048+ 596,    0*2048+ 982,    0*2048+1268,
  24*2048+  70,   27*2048+ 333,    0*2048+ 996,    0*2048+1269,
  20*2048+ 682,    0*2048+ 884,    9*2048+ 907,    0*2048+1270,
  24*2048+ 395,   35*2048+ 471,    0*2048+ 895,    0*2048+1271,
  21*2048+   9,   34*2048+ 645,    0*2048+ 908,    0*2048+1272,
  22*2048+ 533,    0*2048+ 918,   41*2048+ 919,    0*2048+1273,
  14*2048+ 622,    0*2048+ 932,    2*2048+ 983,    0*2048+1274,
  39*2048+ 307,    3*2048+ 920,    0*2048+ 945,    0*2048+1275,
  44*2048+ 134,   12*2048+ 695,    0*2048+ 957,    0*2048+1276,
  26*2048+ 497,   22*2048+ 708,    0*2048+ 971,    0*2048+1277,
  18*2048+ 721,    7*2048+ 958,    0*2048+ 984,    0*2048+1278,
  45*2048+ 195,   15*2048+ 484,    0*2048+ 997,    0*2048+1279,

   0*2048+  14,    0*2048+  30,    0*2048+1392,
   0*2048+  31,    0*2048+  46,    0*2048+1393,
   0*2048+  47,    0*2048+  62,    0*2048+1394,
   0*2048+  63,    0*2048+  81,    0*2048+1395,
   0*2048+  82,    0*2048+  99,    0*2048+1396,
   0*2048+ 100,    0*2048+ 118,    0*2048+1397,
   0*2048+ 119,    0*2048+ 135,    0*2048+1398,
   0*2048+ 136,    0*2048+ 151,    0*2048+1399,
   0*2048+ 152,    0*2048+ 167,    0*2048+1400,
   0*2048+ 168,    0*2048+ 183,    0*2048+1401,
   0*2048+ 184,    0*2048+ 199,    0*2048+1402,
   0*2048+ 200,    0*2048+ 218,    0*2048+1403,
   0*2048+ 219,    0*2048+ 236,    0*2048+1404,
   0*2048+ 237,    0*2048+ 255,    0*2048+1405,
   0*2048+ 256,    0*2048+ 272,    0*2048+1406,
   0*2048+ 273,    0*2048+ 288,    0*2048+1407,
   0*2048+ 289,    0*2048+ 304,    0*2048+1408,
   0*2048+ 305,    0*2048+ 320,    0*2048+1409,
   0*2048+ 321,    0*2048+ 336,    0*2048+1410,
   0*2048+ 337,    0*2048+ 355,    0*2048+1411,
   0*2048+ 356,    0*2048+ 373,    0*2048+1412,
   0*2048+ 374,    0*2048+ 392,    0*2048+1413,
   0*2048+ 393,    0*2048+ 409,    0*2048+1414,
   0*2048+ 410,    0*2048+ 425,    0*2048+1415,
   0*2048+ 426,    0*2048+ 441,    0*2048+1416,
   0*2048+ 442,    0*2048+ 457,    0*2048+1417,
   0*2048+ 458,    0*2048+ 473,    0*2048+1418,
   0*2048+ 474,    0*2048+ 492,    0*2048+1419,
   0*2048+ 493,    0*2048+ 510,    0*2048+1420,
   0*2048+ 511,    0*2048+ 529,    0*2048+1421,
   0*2048+ 530,    0*2048+ 546,    0*2048+1422,
   0*2048+ 547,    0*2048+ 562,    0*2048+1423,
   0*2048+ 563,    0*2048+ 578,    0*2048+1424,
   0*2048+ 579,    0*2048+ 594,    0*2048+1425,
   0*2048+ 595,    0*2048+ 610,    0*2048+1426,
   0*2048+ 611,    0*2048+ 629,    0*2048+1427,
   0*2048+ 630,    0*2048+ 647,    0*2048+1428,
   0*2048+ 648,    0*2048+ 666,    0*2048+1429,
   0*2048+ 667,    0*2048+ 683,    0*2048+1430,
   0*2048+ 684,    0*2048+ 699,    0*2048+1431,
   0*2048+ 700,    0*2048+ 715,    0*2048+1432,
   0*2048+ 716,    0*2048+ 731,    0*2048+1433,
   0*2048+ 732,    0*2048+ 747,    0*2048+1434,
   0*2048+ 748,    0*2048+ 766,    0*2048+1435,
   0*2048+ 767,    0*2048+ 784,    0*2048+1436,
   0*2048+ 785,    0*2048+ 803,    0*2048+1437,
   0*2048+ 804,    0*2048+ 820,    0*2048+1438,
   0*2048+ 821,    0*2048+ 836,    0*2048+1439,
   0*2048+ 837,    0*2048+ 852,    0*2048+1440,
   0*2048+ 853,    0*2048+ 868,    0*2048+1441,
   0*2048+ 869,    0*2048+ 884,    0*2048+1442,
   0*2048+ 885,    0*2048+ 903,    0*2048+1443,
   0*2048+ 904,    0*2048+ 921,    0*2048+1444,
   0*2048+ 922,    0*2048+ 940,    0*2048+1445,
   0*2048+ 941,    0*2048+ 957,    0*2048+1446,
   0*2048+ 958,    0*2048+ 973,    0*2048+1447,
   0*2048+ 974,    0*2048+ 989,    0*2048+1448,
   0*2048+ 990,    0*2048+1005,    0*2048+1449,
   0*2048+1006,    0*2048+1021,    0*2048+1450,
   0*2048+1022,    0*2048+1040,    0*2048+1451,
   0*2048+1041,    0*2048+1058,    0*2048+1452,
   0*2048+1059,    0*2048+1077,    0*2048+1453,
   0*2048+1078,    0*2048+1094,    0*2048+1454,
   1*2048+  15,    0*2048+1095,    0*2048+1455,
   0*2048+  64,   30*2048+ 101,   38*2048+ 257,    0*2048+1097,
   0*2048+  83,   19*2048+ 137,    6*2048+ 512,    0*2048+1098,
  33*2048+  32,    0*2048+ 102,   13*2048+ 169,    0*2048+1099,
   0*2048+ 120,    3*2048+ 338,    8*2048+1042,    0*2048+1100,
   0*2048+   0,   33*2048+   1,   37*2048+ 258,    0*2048+1101,
   0*2048+  16,   36*2048+ 749,   35*2048+ 786,    0*2048+1102,
   0*2048+  33,    8*2048+ 564,   12*2048+ 871,    0*2048+1103,
   0*2048+  49,    2*2048+ 259,   19*2048+ 822,    0*2048+1104,
   0*2048+  65,   35*2048+ 306,   26*2048+ 631,    0*2048+1105,
  15*2048+  66,    0*2048+  84,    2*2048+ 650,    0*2048+1106,
   0*2048+ 103,   37*2048+ 768,    1*2048+ 854,    0*2048+1107,
  35*2048+  50,    0*2048+ 121,    1*2048+ 290,    0*2048+1108,
   0*2048+   2,   19*2048+ 494,   24*2048+ 769,    0*2048+1109,
   0*2048+  17,   12*2048+ 122,    2*2048+ 702,    0*2048+1110,
   0*2048+  34,   17*2048+ 274,   26*2048+ 548,    0*2048+1111,
   0*2048+  51,   44*2048+ 260,   29*2048+ 991,    0*2048+1112,
   0*2048+  67,    8*2048+ 339,   22*2048+ 717,    0*2048+1113,
   0*2048+  85,   15*2048+ 238,    1*2048+ 459,    0*2048+1114,
   0*2048+ 104,    7*2048+ 838,   34*2048+ 886,    0*2048+1115,
   0*2048+ 123,   36*2048+ 375,   24*2048+ 733,    0*2048+1116,
   0*2048+   3,    4*2048+   4,   38*2048+ 855,    0*2048+1117,
   0*2048+  18,   17*2048+ 495,   19*2048+ 770,    0*2048+1118,
   0*2048+  35,   19*2048+ 703,   25*2048+ 992,    0*2048+1119,
   0*2048+  52,   23*2048+ 105,   19*2048+ 154,    0*2048+1120,
   0*2048+  68,   39*2048+ 261,   15*2048+ 340,    0*2048+1121,
   0*2048+  86,   36*2048+ 275,   41*2048+ 872,    0*2048+1122,
   0*2048+ 106,    6*2048+ 873,   19*2048+1060,    0*2048+1123,
   0*2048+ 124,    3*2048+ 612,    7*2048+ 942,    0*2048+1124,
   0*2048+   5,   37*2048+  19,   29*2048+ 496,    0*2048+1125,
   0*2048+  20,    7*2048+ 596,    0*2048+ 975,    0*2048+1126,
   0*2048+  36,   13*2048+ 107,   16*2048+ 443,    0*2048+1127,
   0*2048+  53,   31*2048+ 108,   19*2048+ 262,    0*2048+1128,
   0*2048+  69,    1*2048+  70,   27*2048+ 170,    0*2048+1129,
   0*2048+  87,   37*2048+ 412,   14*2048+ 943,    0*2048+1130,
  10*2048+  88,    0*2048+ 109,    2*2048+ 597,    0*2048+1131,
   0*2048+ 125,   41*2048+ 341,   26*2048+ 685,    0*2048+1132,
   0*2048+ 204,   30*2048+ 239,   38*2048+ 394,    0*2048+1134,
   0*2048+ 221,   19*2048+ 276,    6*2048+ 651,    0*2048+1135,
  33*2048+ 171,    0*2048+ 240,   13*2048+ 307,    0*2048+1136,
   9*2048+  89,    0*2048+ 263,    3*2048+ 475,    0*2048+1137,
   0*2048+ 138,   33*2048+ 139,   37*2048+ 395,    0*2048+1138,
   0*2048+ 155,   36*2048+ 887,   35*2048+ 924,    0*2048+1139,
   0*2048+ 172,    8*2048+ 704,   12*2048+1008,    0*2048+1140,
   0*2048+ 186,    2*2048+ 396,   19*2048+ 959,    0*2048+1141,
   0*2048+ 205,   35*2048+ 444,   26*2048+ 771,    0*2048+1142,
  15*2048+ 206,    0*2048+ 222,    2*2048+ 788,    0*2048+1143,
   0*2048+ 241,   37*2048+ 906,    1*2048+ 993,    0*2048+1144,
  35*2048+ 187,    0*2048+ 264,    1*2048+ 427,    0*2048+1145,
   0*2048+ 140,   19*2048+ 632,   24*2048+ 907,    0*2048+1146,
   0*2048+ 156,   12*2048+ 265,    2*2048+ 840,    0*2048+1147,
   0*2048+ 173,   17*2048+ 413,   26*2048+ 686,    0*2048+1148,
  30*2048+  37,    0*2048+ 188,   44*2048+ 397,    0*2048+1149,
   0*2048+ 207,    8*2048+ 476,   22*2048+ 856,    0*2048+1150,
   0*2048+ 223,   15*2048+ 376,    1*2048+ 598,    0*2048+1151,
   0*2048+ 242,    7*2048+ 976,   34*2048+1023,    0*2048+1152,
   0*2048+ 266,   36*2048+ 513,   24*2048+ 874,    0*2048+1153,
   0*2048+ 141,    4*2048+ 142,   38*2048+ 994,    0*2048+1154,
   0*2048+ 157,   17*2048+ 633,   19*2048+ 908,    0*2048+1155,
  26*2048+  38,    0*2048+ 174,   19*2048+ 841,    0*2048+1156,
   0*2048+ 189,   23*2048+ 243,   19*2048+ 292,    0*2048+1157,
   0*2048+ 208,   39*2048+ 398,   15*2048+ 477,    0*2048+1158,
   0*2048+ 224,   36*2048+ 414,   41*2048+1009,    0*2048+1159,
  20*2048+ 110,    0*2048+ 244,    6*2048+1010,    0*2048+1160,
   0*2048+ 267,    3*2048+ 750,    7*2048+1079,    0*2048+1161,
   0*2048+ 143,   37*2048+ 158,   29*2048+ 634,    0*2048+1162,
   1*2048+  21,    0*2048+ 159,    7*2048+ 734,    0*2048+1163,
   0*2048+ 175,   13*2048+ 245,   16*2048+ 580,    0*2048+1164,
   0*2048+ 190,   31*2048+ 246,   19*2048+ 399,    0*2048+1165,
   0*2048+ 209,    1*2048+ 210,   27*2048+ 308,    0*2048+1166,
   0*2048+ 225,   37*2048+ 550,   14*2048+1080,    0*2048+1167,
  10*2048+ 226,    0*2048+ 247,    2*2048+ 735,    0*2048+1168,
   0*2048+ 268,   41*2048+ 478,   26*2048+ 823,    0*2048+1169,
   0*2048+ 345,   30*2048+ 377,   38*2048+ 531,    0*2048+1171,
   0*2048+ 358,   19*2048+ 415,    6*2048+ 789,    0*2048+1172,
  33*2048+ 309,    0*2048+ 378,   13*2048+ 445,    0*2048+1173,
   9*2048+ 227,    0*2048+ 400,    3*2048+ 613,    0*2048+1174,
   0*2048+ 277,   33*2048+ 278,   37*2048+ 532,    0*2048+1175,
   0*2048+ 293,   36*2048+1024,   35*2048+1062,    0*2048+1176,
  13*2048+  55,    0*2048+ 310,    8*2048+ 842,    0*2048+1177,
  20*2048+   6,    0*2048+ 323,    2*2048+ 533,    0*2048+1178,
   0*2048+ 346,   35*2048+ 581,   26*2048+ 909,    0*2048+1179,
  15*2048+ 347,    0*2048+ 359,    2*2048+ 926,    0*2048+1180,
   2*2048+  39,    0*2048+ 379,   37*2048+1044,    0*2048+1181,
  35*2048+ 324,    0*2048+ 401,    1*2048+ 565,    0*2048+1182,
   0*2048+ 279,   19*2048+ 772,   24*2048+1045,    0*2048+1183,
   0*2048+ 294,   12*2048+ 402,    2*2048+ 978,    0*2048+1184,
   0*2048+ 311,   17*2048+ 551,   26*2048+ 824,    0*2048+1185,
  30*2048+ 176,    0*2048+ 325,   44*2048+ 534,    0*2048+1186,
   0*2048+ 348,    8*2048+ 614,   22*2048+ 995,    0*2048+1187,
   0*2048+ 360,   15*2048+ 514,    1*2048+ 736,    0*2048+1188,
   8*2048+  22,   35*2048+  71,    0*2048+ 380,    0*2048+1189,
   0*2048+ 403,   36*2048+ 652,   24*2048+1011,    0*2048+1190,
  39*2048+  40,    0*2048+ 280,    4*2048+ 281,    0*2048+1191,
   0*2048+ 295,   17*2048+ 773,   19*2048+1046,    0*2048+1192,
  26*2048+ 177,    0*2048+ 312,   19*2048+ 979,    0*2048+1193,
   0*2048+ 326,   23*2048+ 381,   19*2048+ 429,    0*2048+1194,
   0*2048+ 349,   39*2048+ 535,   15*2048+ 615,    0*2048+1195,
  42*2048+  56,    0*2048+ 361,   36*2048+ 552,    0*2048+1196,
   7*2048+  57,   20*2048+ 248,    0*2048+ 382,    0*2048+1197,
   8*2048+ 126,    0*2048+ 404,    3*2048+ 888,    0*2048+1198,
   0*2048+ 282,   37*2048+ 296,   29*2048+ 774,    0*2048+1199,
   1*2048+ 160,    0*2048+ 297,    7*2048+ 875,    0*2048+1200,
   0*2048+ 313,   13*2048+ 383,   16*2048+ 718,    0*2048+1201,
   0*2048+ 327,   31*2048+ 384,   19*2048+ 536,    0*2048+1202,
   0*2048+ 350,    1*2048+ 351,   27*2048+ 446,    0*2048+1203,
  15*2048+ 127,    0*2048+ 362,   37*2048+ 688,    0*2048+1204,
  10*2048+ 363,    0*2048+ 385,    2*2048+ 876,    0*2048+1205,
   0*2048+ 405,   41*2048+ 616,   26*2048+ 960,    0*2048+1206,
   0*2048+ 482,   30*2048+ 515,   38*2048+ 668,    0*2048+1208,
   0*2048+ 498,   19*2048+ 553,    6*2048+ 927,    0*2048+1209,
  33*2048+ 447,    0*2048+ 516,   13*2048+ 582,    0*2048+1210,
   9*2048+ 364,    0*2048+ 537,    3*2048+ 751,    0*2048+1211,
   0*2048+ 416,   33*2048+ 417,   37*2048+ 669,    0*2048+1212,
  37*2048+  72,   36*2048+ 112,    0*2048+ 430,    0*2048+1213,
  13*2048+ 192,    0*2048+ 448,    8*2048+ 980,    0*2048+1214,
  20*2048+ 144,    0*2048+ 461,    2*2048+ 670,    0*2048+1215,
   0*2048+ 483,   35*2048+ 719,   26*2048+1047,    0*2048+1216,
  15*2048+ 484,    0*2048+ 499,    2*2048+1064,    0*2048+1217,
  38*2048+  91,    2*2048+ 178,    0*2048+ 517,    0*2048+1218,
  35*2048+ 462,    0*2048+ 538,    1*2048+ 705,    0*2048+1219,
  25*2048+  92,    0*2048+ 418,   19*2048+ 910,    0*2048+1220,
   3*2048+  24,    0*2048+ 431,   12*2048+ 539,    0*2048+1221,
   0*2048+ 449,   17*2048+ 689,   26*2048+ 961,    0*2048+1222,
  30*2048+ 314,    0*2048+ 463,   44*2048+ 671,    0*2048+1223,
  23*2048+  41,    0*2048+ 485,    8*2048+ 752,    0*2048+1224,
   0*2048+ 500,   15*2048+ 653,    1*2048+ 877,    0*2048+1225,
   8*2048+ 161,   35*2048+ 211,    0*2048+ 518,    0*2048+1226,
  25*2048+  58,    0*2048+ 540,   36*2048+ 790,    0*2048+1227,
  39*2048+ 179,    0*2048+ 419,    4*2048+ 420,    0*2048+1228,
  20*2048+  93,    0*2048+ 432,   17*2048+ 911,    0*2048+1229,
  20*2048+  25,   26*2048+ 315,    0*2048+ 450,    0*2048+1230,
   0*2048+ 464,   23*2048+ 519,   19*2048+ 567,    0*2048+1231,
   0*2048+ 486,   39*2048+ 672,   15*2048+ 753,    0*2048+1232,
  42*2048+ 193,    0*2048+ 501,   36*2048+ 690,    0*2048+1233,
   7*2048+ 194,   20*2048+ 386,    0*2048+ 520,    0*2048+1234,
   8*2048+ 269,    0*2048+ 541,    3*2048+1025,    0*2048+1235,
   0*2048+ 421,   37*2048+ 433,   29*2048+ 912,    0*2048+1236,
   1*2048+ 298,    0*2048+ 434,    7*2048+1012,    0*2048+1237,
   0*2048+ 451,   13*2048+ 521,   16*2048+ 857,    0*2048+1238,
   0*2048+ 465,   31*2048+ 522,   19*2048+ 673,    0*2048+1239,
   0*2048+ 487,    1*2048+ 488,   27*2048+ 583,    0*2048+1240,
  15*2048+ 270,    0*2048+ 502,   37*2048+ 826,    0*2048+1241,
  10*2048+ 503,    0*2048+ 523,    2*2048+1013,    0*2048+1242,
  27*2048+   7,    0*2048+ 542,   41*2048+ 754,    0*2048+1243,
   0*2048+ 620,   30*2048+ 654,   38*2048+ 806,    0*2048+1245,
   0*2048+ 636,   19*2048+ 691,    6*2048+1065,    0*2048+1246,
  33*2048+ 584,    0*2048+ 655,   13*2048+ 720,    0*2048+1247,
   9*2048+ 504,    0*2048+ 674,    3*2048+ 889,    0*2048+1248,
   0*2048+ 554,   33*2048+ 555,   37*2048+ 807,    0*2048+1249,
  37*2048+ 212,   36*2048+ 250,    0*2048+ 568,    0*2048+1250,
   9*2048+  26,   13*2048+ 329,    0*2048+ 585,    0*2048+1251,
  20*2048+ 283,    0*2048+ 600,    2*2048+ 808,    0*2048+1252,
  27*2048+  94,    0*2048+ 621,   35*2048+ 858,    0*2048+1253,
   3*2048+ 114,   15*2048+ 622,    0*2048+ 637,    0*2048+1254,
  38*2048+ 229,    2*2048+ 316,    0*2048+ 656,    0*2048+1255,
  35*2048+ 601,    0*2048+ 675,    1*2048+ 843,    0*2048+1256,
  25*2048+ 230,    0*2048+ 556,   19*2048+1048,    0*2048+1257,
   3*2048+ 163,    0*2048+ 569,   12*2048+ 676,    0*2048+1258,
  27*2048+   8,    0*2048+ 586,   17*2048+ 827,    0*2048+1259,
  30*2048+ 452,    0*2048+ 602,   44*2048+ 809,    0*2048+1260,
  23*2048+ 180,    0*2048+ 623,    8*2048+ 890,    0*2048+1261,
   0*2048+ 638,   15*2048+ 791,    1*2048+1014,    0*2048+1262,
   8*2048+ 299,   35*2048+ 352,    0*2048+ 657,    0*2048+1263,
  25*2048+ 195,    0*2048+ 677,   36*2048+ 928,    0*2048+1264,
  39*2048+ 317,    0*2048+ 557,    4*2048+ 558,    0*2048+1265,
  20*2048+ 231,    0*2048+ 570,   17*2048+1049,    0*2048+1266,
  20*2048+ 164,   26*2048+ 453,    0*2048+ 587,    0*2048+1267,
   0*2048+ 603,   23*2048+ 658,   19*2048+ 707,    0*2048+1268,
   0*2048+ 624,   39*2048+ 810,   15*2048+ 891,    0*2048+1269,
  42*2048+ 330,    0*2048+ 639,   36*2048+ 828,    0*2048+1270,
   7*2048+ 331,   20*2048+ 524,    0*2048+ 659,    0*2048+1271,
   4*2048+  73,    8*2048+ 406,    0*2048+ 678,    0*2048+1272,
   0*2048+ 559,   37*2048+ 571,   29*2048+1050,    0*2048+1273,
   8*2048+  59,    1*2048+ 435,    0*2048+ 572,    0*2048+1274,
   0*2048+ 588,   13*2048+ 660,   16*2048+ 996,    0*2048+1275,
   0*2048+ 604,   31*2048+ 661,   19*2048+ 811,    0*2048+1276,
   0*2048+ 625,    1*2048+ 626,   27*2048+ 721,    0*2048+1277,
  15*2048+ 407,    0*2048+ 640,   37*2048+ 963,    0*2048+1278,
   3*2048+  60,   10*2048+ 641,    0*2048+ 662,    0*2048+1279,
  27*2048+ 145,    0*2048+ 679,   41*2048+ 892,    0*2048+1280,
   0*2048+ 758,   30*2048+ 792,   38*2048+ 945,    0*2048+1282,
   7*2048+ 115,    0*2048+ 776,   19*2048+ 829,    0*2048+1283,
  33*2048+ 722,    0*2048+ 793,   13*2048+ 859,    0*2048+1284,
   9*2048+ 642,    0*2048+ 812,    3*2048+1026,    0*2048+1285,
   0*2048+ 692,   33*2048+ 693,   37*2048+ 946,    0*2048+1286,
  37*2048+ 353,   36*2048+ 388,    0*2048+ 708,    0*2048+1287,
   9*2048+ 165,   13*2048+ 467,    0*2048+ 723,    0*2048+1288,
  20*2048+ 422,    0*2048+ 738,    2*2048+ 947,    0*2048+1289,
  27*2048+ 232,    0*2048+ 759,   35*2048+ 997,    0*2048+1290,
   3*2048+ 252,   15*2048+ 760,    0*2048+ 777,    0*2048+1291,
  38*2048+ 366,    2*2048+ 454,    0*2048+ 794,    0*2048+1292,
  35*2048+ 739,    0*2048+ 813,    1*2048+ 981,    0*2048+1293,
  20*2048+  95,   25*2048+ 367,    0*2048+ 694,    0*2048+1294,
   3*2048+ 301,    0*2048+ 709,   12*2048+ 814,    0*2048+1295,
  27*2048+ 146,    0*2048+ 724,   17*2048+ 964,    0*2048+1296,
  30*2048+ 589,    0*2048+ 740,   44*2048+ 948,    0*2048+1297,
  23*2048+ 318,    0*2048+ 761,    8*2048+1027,    0*2048+1298,
   2*2048+  61,    0*2048+ 778,   15*2048+ 929,    0*2048+1299,
   8*2048+ 436,   35*2048+ 489,    0*2048+ 795,    0*2048+1300,
  25*2048+ 332,    0*2048+ 815,   36*2048+1066,    0*2048+1301,
  39*2048+ 455,    0*2048+ 695,    4*2048+ 696,    0*2048+1302,
  18*2048+  96,   20*2048+ 368,    0*2048+ 710,    0*2048+1303,
  20*2048+ 302,   26*2048+ 590,    0*2048+ 725,    0*2048+1304,
   0*2048+ 741,   23*2048+ 796,   19*2048+ 845,    0*2048+1305,
   0*2048+ 762,   39*2048+ 949,   15*2048+1028,    0*2048+1306,
  42*2048+ 468,    0*2048+ 779,   36*2048+ 965,    0*2048+1307,
   7*2048+ 469,   20*2048+ 663,    0*2048+ 797,    0*2048+1308,
   4*2048+ 213,    8*2048+ 543,    0*2048+ 816,    0*2048+1309,
  30*2048+  97,    0*2048+ 697,   37*2048+ 711,    0*2048+1310,
   8*2048+ 196,    1*2048+ 573,    0*2048+ 712,    0*2048+1311,
  17*2048+  42,    0*2048+ 726,   13*2048+ 798,    0*2048+1312,
   0*2048+ 742,   31*2048+ 799,   19*2048+ 950,    0*2048+1313,
   0*2048+ 763,    1*2048+ 764,   27*2048+ 860,    0*2048+1314,
  38*2048+  10,   15*2048+ 544,    0*2048+ 780,    0*2048+1315,
   3*2048+ 197,   10*2048+ 781,    0*2048+ 800,    0*2048+1316,
  27*2048+ 284,    0*2048+ 817,   41*2048+1029,    0*2048+1317,
   0*2048+ 896,   30*2048+ 930,   38*2048+1082,    0*2048+1319,
   7*2048+ 253,    0*2048+ 914,   19*2048+ 966,    0*2048+1320,
  33*2048+ 861,    0*2048+ 931,   13*2048+ 998,    0*2048+1321,
   4*2048+  74,    9*2048+ 782,    0*2048+ 951,    0*2048+1322,
   0*2048+ 830,   33*2048+ 831,   37*2048+1083,    0*2048+1323,
  37*2048+ 490,   36*2048+ 526,    0*2048+ 846,    0*2048+1324,
   9*2048+ 303,   13*2048+ 606,    0*2048+ 862,    0*2048+1325,
  20*2048+ 560,    0*2048+ 879,    2*2048+1084,    0*2048+1326,
  36*2048+  43,   27*2048+ 369,    0*2048+ 897,    0*2048+1327,
   3*2048+ 390,   15*2048+ 898,    0*2048+ 915,    0*2048+1328,
  38*2048+ 506,    2*2048+ 591,    0*2048+ 932,    0*2048+1329,
   2*2048+  27,   35*2048+ 880,    0*2048+ 952,    0*2048+1330,
  20*2048+ 233,   25*2048+ 507,    0*2048+ 832,    0*2048+1331,
   3*2048+ 438,    0*2048+ 847,   12*2048+ 953,    0*2048+1332,
  18*2048+  11,   27*2048+ 285,    0*2048+ 863,    0*2048+1333,
  30*2048+ 727,    0*2048+ 881,   44*2048+1085,    0*2048+1334,
   9*2048+  75,   23*2048+ 456,    0*2048+ 899,    0*2048+1335,
   2*2048+ 198,    0*2048+ 916,   15*2048+1067,    0*2048+1336,
   8*2048+ 574,   35*2048+ 627,    0*2048+ 933,    0*2048+1337,
  37*2048+ 116,   25*2048+ 470,    0*2048+ 954,    0*2048+1338,
  39*2048+ 592,    0*2048+ 833,    4*2048+ 834,    0*2048+1339,
  18*2048+ 234,   20*2048+ 508,    0*2048+ 848,    0*2048+1340,
  20*2048+ 439,   26*2048+ 728,    0*2048+ 864,    0*2048+1341,
   0*2048+ 882,   23*2048+ 934,   19*2048+ 983,    0*2048+1342,
  16*2048+  76,    0*2048+ 900,   39*2048+1086,    0*2048+1343,
  37*2048+  12,   42*2048+ 607,    0*2048+ 917,    0*2048+1344,
   7*2048+ 608,   20*2048+ 801,    0*2048+ 935,    0*2048+1345,
   4*2048+ 354,    8*2048+ 680,    0*2048+ 955,    0*2048+1346,
  30*2048+ 235,    0*2048+ 835,   37*2048+ 849,    0*2048+1347,
   8*2048+ 333,    1*2048+ 713,    0*2048+ 850,    0*2048+1348,
  17*2048+ 181,    0*2048+ 865,   13*2048+ 936,    0*2048+1349,
   0*2048+ 883,   31*2048+ 937,   19*2048+1087,    0*2048+1350,
   0*2048+ 901,    1*2048+ 902,   27*2048+ 999,    0*2048+1351,
  38*2048+ 148,   15*2048+ 681,    0*2048+ 918,    0*2048+1352,
   3*2048+ 334,   10*2048+ 919,    0*2048+ 938,    0*2048+1353,
  42*2048+  77,   27*2048+ 423,    0*2048+ 956,    0*2048+1354,
  39*2048+ 129,    0*2048+1033,   30*2048+1068,    0*2048+1356,
  20*2048+  13,    7*2048+ 391,    0*2048+1052,    0*2048+1357,
  14*2048+  44,   33*2048+1000,    0*2048+1069,    0*2048+1358,
   4*2048+ 214,    9*2048+ 920,    0*2048+1088,    0*2048+1359,
  38*2048+ 130,    0*2048+ 967,   33*2048+ 968,    0*2048+1360,
  37*2048+ 628,   36*2048+ 665,    0*2048+ 984,    0*2048+1361,
   9*2048+ 440,   13*2048+ 744,    0*2048+1001,    0*2048+1362,
   3*2048+ 131,   20*2048+ 698,    0*2048+1016,    0*2048+1363,
  36*2048+ 182,   27*2048+ 509,    0*2048+1034,    0*2048+1364,
   3*2048+ 528,   15*2048+1035,    0*2048+1053,    0*2048+1365,
  38*2048+ 644,    2*2048+ 729,    0*2048+1070,    0*2048+1366,
   2*2048+ 166,   35*2048+1017,    0*2048+1089,    0*2048+1367,
  20*2048+ 370,   25*2048+ 645,    0*2048+ 969,    0*2048+1368,
   3*2048+ 576,    0*2048+ 985,   12*2048+1090,    0*2048+1369,
  18*2048+ 149,   27*2048+ 424,    0*2048+1002,    0*2048+1370,
  45*2048+ 132,   30*2048+ 866,    0*2048+1018,    0*2048+1371,
   9*2048+ 215,   23*2048+ 593,    0*2048+1036,    0*2048+1372,
  16*2048+ 117,    2*2048+ 335,    0*2048+1054,    0*2048+1373,
   8*2048+ 714,   35*2048+ 765,    0*2048+1071,    0*2048+1374,
  37*2048+ 254,   25*2048+ 609,    0*2048+1091,    0*2048+1375,
  39*2048+ 730,    0*2048+ 970,    4*2048+ 971,    0*2048+1376,
  18*2048+ 371,   20*2048+ 646,    0*2048+ 986,    0*2048+1377,
  20*2048+ 577,   26*2048+ 867,    0*2048+1003,    0*2048+1378,
  20*2048+  29,    0*2048+1019,   23*2048+1072,    0*2048+1379,
  40*2048+ 133,   16*2048+ 216,    0*2048+1037,    0*2048+1380,
  37*2048+ 150,   42*2048+ 745,    0*2048+1055,    0*2048+1381,
   7*2048+ 746,   20*2048+ 939,    0*2048+1073,    0*2048+1382,
   4*2048+ 491,    8*2048+ 818,    0*2048+1092,    0*2048+1383,
  30*2048+ 372,    0*2048+ 972,   37*2048+ 987,    0*2048+1384,
   8*2048+ 471,    1*2048+ 851,    0*2048+ 988,    0*2048+1385,
  17*2048+ 319,    0*2048+1004,   13*2048+1074,    0*2048+1386,
  20*2048+ 134,    0*2048+1020,   31*2048+1075,    0*2048+1387,
  28*2048+  45,    0*2048+1038,    1*2048+1039,    0*2048+1388,
  38*2048+ 287,   15*2048+ 819,    0*2048+1056,    0*2048+1389,
   3*2048+ 472,   10*2048+1057,    0*2048+1076,    0*2048+1390,
  42*2048+ 217,   27*2048+ 561,    0*2048+1093,    0*2048+1391,
   0*2048+  48,   23*2048+ 153,   14*2048+ 201,   11*2048+ 202,   39*2048+ 203,    5*2048+ 220,   35*2048+ 411,   26*2048+ 649,   37*2048+ 701,    8*2048+ 805,    7*2048+ 870,   43*2048+ 905,   19*2048+ 923,    0*2048+1096,
   0*2048+ 185,   23*2048+ 291,   14*2048+ 342,   11*2048+ 343,   39*2048+ 344,    5*2048+ 357,   35*2048+ 549,   26*2048+ 787,   37*2048+ 839,    8*2048+ 944,    7*2048+1007,   43*2048+1043,   19*2048+1061,    0*2048+1133,
   8*2048+  54,   44*2048+  90,   20*2048+ 111,    0*2048+ 322,   23*2048+ 428,   14*2048+ 479,   11*2048+ 480,   39*2048+ 481,    5*2048+ 497,   35*2048+ 687,   26*2048+ 925,   37*2048+ 977,    8*2048+1081,    0*2048+1170,
  38*2048+  23,    9*2048+ 128,    8*2048+ 191,   44*2048+ 228,   20*2048+ 249,    0*2048+ 460,   23*2048+ 566,   14*2048+ 617,   11*2048+ 618,   39*2048+ 619,    5*2048+ 635,   35*2048+ 825,   26*2048+1063,    0*2048+1207,
  27*2048+ 113,   38*2048+ 162,    9*2048+ 271,    8*2048+ 328,   44*2048+ 365,   20*2048+ 387,    0*2048+ 599,   23*2048+ 706,   14*2048+ 755,   11*2048+ 756,   39*2048+ 757,    5*2048+ 775,   35*2048+ 962,    0*2048+1244,
  36*2048+   9,   27*2048+ 251,   38*2048+ 300,    9*2048+ 408,    8*2048+ 466,   44*2048+ 505,   20*2048+ 525,    0*2048+ 737,   23*2048+ 844,   14*2048+ 893,   11*2048+ 894,   39*2048+ 895,    5*2048+ 913,    0*2048+1281,
  36*2048+ 147,   27*2048+ 389,   38*2048+ 437,    9*2048+ 545,    8*2048+ 605,   44*2048+ 643,   20*2048+ 664,    0*2048+ 878,   23*2048+ 982,   14*2048+1030,   11*2048+1031,   39*2048+1032,    5*2048+1051,    0*2048+1318,
  24*2048+  28,   15*2048+  78,   12*2048+  79,   40*2048+  80,    6*2048+  98,   36*2048+ 286,   27*2048+ 527,   38*2048+ 575,    9*2048+ 682,    8*2048+ 743,   44*2048+ 783,   20*2048+ 802,    0*2048+1015,    0*2048+1355,

   0*2048+  25,    0*2048+  52,    0*2048+1400,
   0*2048+  53,    0*2048+  79,    0*2048+1401,
   0*2048+  80,    0*2048+ 106,    0*2048+1402,
   0*2048+ 107,    0*2048+ 133,    0*2048+1403,
   0*2048+ 134,    0*2048+ 160,    0*2048+1404,
   0*2048+ 161,    0*2048+ 187,    0*2048+1405,
   0*2048+ 188,    0*2048+ 214,    0*2048+1406,
   0*2048+ 215,    0*2048+ 241,    0*2048+1407,
   0*2048+ 242,    0*2048+ 268,    0*2048+1408,
   0*2048+ 269,    0*2048+ 295,    0*2048+1409,
   0*2048+ 296,    0*2048+ 322,    0*2048+1410,
   0*2048+ 323,    0*2048+ 349,    0*2048+1411,
   0*2048+ 350,    0*2048+ 376,    0*2048+1412,
   0*2048+ 377,    0*2048+ 403,    0*2048+1413,
   0*2048+ 404,    0*2048+ 430,    0*2048+1414,
   0*2048+ 431,    0*2048+ 457,    0*2048+1415,
   0*2048+ 458,    0*2048+ 484,    0*2048+1416,
   0*2048+ 485,    0*2048+ 511,    0*2048+1417,
   0*2048+ 512,    0*2048+ 538,    0*2048+1418,
   0*2048+ 539,    0*2048+ 565,    0*2048+1419,
   0*2048+ 566,    0*2048+ 592,    0*2048+1420,
   0*2048+ 593,    0*2048+ 619,    0*2048+1421,
   0*2048+ 620,    0*2048+ 646,    0*2048+1422,
   0*2048+ 647,    0*2048+ 673,    0*2048+1423,
   0*2048+ 674,    0*2048+ 700,    0*2048+1424,
   0*2048+ 701,    0*2048+ 727,    0*2048+1425,
   0*2048+ 728,    0*2048+ 754,    0*2048+1426,
   0*2048+ 755,    0*2048+ 781,    0*2048+1427,
   0*2048+ 782,    0*2048+ 808,    0*2048+1428,
   0*2048+ 809,    0*2048+ 835,    0*2048+1429,
   0*2048+ 836,    0*2048+ 862,    0*2048+1430,
   0*2048+ 863,    0*2048+ 889,    0*2048+1431,
   0*2048+ 890,    0*2048+ 916,    0*2048+1432,
   0*2048+ 917,    0*2048+ 943,    0*2048+1433,
   0*2048+ 944,    0*2048+ 970,    0*2048+1434,
   0*2048+ 971,    0*2048+ 997,    0*2048+1435,
   0*2048+ 998,    0*2048+1024,    0*2048+1436,
   0*2048+1025,    0*2048+1051,    0*2048+1437,
   0*2048+1052,    0*2048+1078,    0*2048+1438,
   1*2048+  26,    0*2048+1079,    0*2048+1439,
   0*2048+   1,   23*2048+ 164,   39*2048+ 486,    0*2048+1085,
   0*2048+  28,   34*2048+ 379,   19*2048+ 460,    0*2048+1086,
   0*2048+  56,   15*2048+ 216,    3*2048+ 837,    0*2048+1087,
   0*2048+  83,    5*2048+ 271,   29*2048+ 945,    0*2048+1088,
   0*2048+ 109,   37*2048+ 110,   17*2048+ 324,    0*2048+1089,
   0*2048+   2,   12*2048+ 217,   10*2048+ 729,    0*2048+1090,
   0*2048+  29,   28*2048+ 111,   20*2048+ 756,    0*2048+1091,
   0*2048+  57,   34*2048+ 165,   21*2048+ 918,    0*2048+1092,
   0*2048+  84,   37*2048+ 540,   20*2048+ 946,    0*2048+1093,
   0*2048+ 112,   37*2048+ 432,   12*2048+ 594,    0*2048+1094,
   0*2048+   3,   25*2048+ 166,   42*2048+ 568,    0*2048+1095,
   0*2048+  30,    2*2048+ 461,   28*2048+ 947,    0*2048+1096,
   0*2048+  58,   35*2048+  85,   16*2048+ 462,    0*2048+1097,
   0*2048+  86,   36*2048+ 351,   15*2048+ 649,    0*2048+1098,
   0*2048+ 113,   37*2048+ 405,   10*2048+ 783,    0*2048+1099,
   0*2048+   4,   20*2048+ 244,    9*2048+ 675,    0*2048+1100,
   0*2048+  31,    9*2048+ 189,    3*2048+ 838,    0*2048+1101,
   0*2048+  59,    5*2048+  60,   33*2048+  87,    0*2048+1102,
  24*2048+   5,    0*2048+  88,    7*2048+1027,    0*2048+1103,
   0*2048+ 114,   36*2048+ 297,   25*2048+1053,    0*2048+1104,
   0*2048+   6,   43*2048+  61,   27*2048+ 487,    0*2048+1105,
   0*2048+  32,   25*2048+ 406,   35*2048+ 757,    0*2048+1106,
   0*2048+  62,   39*2048+ 115,   31*2048+ 569,    0*2048+1107,
   0*2048+  89,   13*2048+ 650,   29*2048+ 810,    0*2048+1108,
   0*2048+ 116,   31*2048+ 167,   36*2048+ 865,    0*2048+1109,
   0*2048+   7,   12*2048+ 758,   15*2048+ 811,    0*2048+1110,
   0*2048+  33,   10*2048+ 570,   42*2048+ 651,    0*2048+1111,
   0*2048+  63,    7*2048+ 117,   22*2048+ 488,    0*2048+1112,
   0*2048+  90,   14*2048+ 463,    9*2048+ 866,    0*2048+1113,
   0*2048+ 118,   28*2048+ 948,   13*2048+ 972,    0*2048+1114,
   0*2048+   8,   25*2048+   9,   15*2048+ 839,    0*2048+1115,
   0*2048+  34,   34*2048+ 218,   18*2048+ 325,    0*2048+1116,
   0*2048+  64,   33*2048+ 219,    8*2048+ 245,    0*2048+1117,
   0*2048+  91,   12*2048+ 702,   37*2048+ 949,    0*2048+1118,
   0*2048+ 119,   29*2048+ 326,   27*2048+ 652,    0*2048+1119,
   0*2048+ 138,   23*2048+ 300,   39*2048+ 621,    0*2048+1125,
   0*2048+ 169,   34*2048+ 514,   19*2048+ 596,    0*2048+1126,
   0*2048+ 192,   15*2048+ 352,    3*2048+ 973,    0*2048+1127,
  30*2048+  10,    0*2048+ 222,    5*2048+ 408,    0*2048+1128,
   0*2048+ 247,   37*2048+ 248,   17*2048+ 464,    0*2048+1129,
   0*2048+ 139,   12*2048+ 353,   10*2048+ 867,    0*2048+1130,
   0*2048+ 170,   28*2048+ 249,   20*2048+ 892,    0*2048+1131,
   0*2048+ 193,   34*2048+ 301,   21*2048+1054,    0*2048+1132,
  21*2048+  11,    0*2048+ 223,   37*2048+ 676,    0*2048+1133,
   0*2048+ 250,   37*2048+ 571,   12*2048+ 730,    0*2048+1134,
   0*2048+ 140,   25*2048+ 302,   42*2048+ 704,    0*2048+1135,
  29*2048+  12,    0*2048+ 171,    2*2048+ 597,    0*2048+1136,
   0*2048+ 194,   35*2048+ 224,   16*2048+ 598,    0*2048+1137,
   0*2048+ 225,   36*2048+ 489,   15*2048+ 785,    0*2048+1138,
   0*2048+ 251,   37*2048+ 541,   10*2048+ 919,    0*2048+1139,
   0*2048+ 141,   20*2048+ 381,    9*2048+ 812,    0*2048+1140,
   0*2048+ 172,    9*2048+ 327,    3*2048+ 974,    0*2048+1141,
   0*2048+ 195,    5*2048+ 196,   33*2048+ 226,    0*2048+1142,
   8*2048+  93,   24*2048+ 142,    0*2048+ 227,    0*2048+1143,
  26*2048+ 120,    0*2048+ 252,   36*2048+ 433,    0*2048+1144,
   0*2048+ 143,   43*2048+ 197,   27*2048+ 622,    0*2048+1145,
   0*2048+ 173,   25*2048+ 542,   35*2048+ 893,    0*2048+1146,
   0*2048+ 198,   39*2048+ 253,   31*2048+ 705,    0*2048+1147,
   0*2048+ 228,   13*2048+ 786,   29*2048+ 950,    0*2048+1148,
   0*2048+ 254,   31*2048+ 303,   36*2048+1000,    0*2048+1149,
   0*2048+ 144,   12*2048+ 894,   15*2048+ 951,    0*2048+1150,
   0*2048+ 174,   10*2048+ 706,   42*2048+ 787,    0*2048+1151,
   0*2048+ 199,    7*2048+ 255,   22*2048+ 623,    0*2048+1152,
   0*2048+ 229,   14*2048+ 599,    9*2048+1001,    0*2048+1153,
  29*2048+  13,   14*2048+  35,    0*2048+ 256,    0*2048+1154,
   0*2048+ 145,   25*2048+ 146,   15*2048+ 975,    0*2048+1155,
   0*2048+ 175,   34*2048+ 354,   18*2048+ 465,    0*2048+1156,
   0*2048+ 200,   33*2048+ 355,    8*2048+ 382,    0*2048+1157,
  38*2048+  14,    0*2048+ 230,   12*2048+ 840,    0*2048+1158,
   0*2048+ 257,   29*2048+ 466,   27*2048+ 788,    0*2048+1159,
   0*2048+ 275,   23*2048+ 436,   39*2048+ 759,    0*2048+1165,
   0*2048+ 305,   34*2048+ 654,   19*2048+ 732,    0*2048+1166,
   4*2048+  36,    0*2048+ 330,   15*2048+ 490,    0*2048+1167,
  30*2048+ 147,    0*2048+ 358,    5*2048+ 544,    0*2048+1168,
   0*2048+ 384,   37*2048+ 385,   17*2048+ 600,    0*2048+1169,
   0*2048+ 276,   12*2048+ 491,   10*2048+1002,    0*2048+1170,
   0*2048+ 306,   28*2048+ 386,   20*2048+1029,    0*2048+1171,
  22*2048+ 121,    0*2048+ 331,   34*2048+ 437,    0*2048+1172,
  21*2048+ 148,    0*2048+ 359,   37*2048+ 813,    0*2048+1173,
   0*2048+ 387,   37*2048+ 707,   12*2048+ 868,    0*2048+1174,
   0*2048+ 277,   25*2048+ 438,   42*2048+ 842,    0*2048+1175,
  29*2048+ 149,    0*2048+ 307,    2*2048+ 733,    0*2048+1176,
   0*2048+ 332,   35*2048+ 360,   16*2048+ 734,    0*2048+1177,
   0*2048+ 361,   36*2048+ 624,   15*2048+ 921,    0*2048+1178,
   0*2048+ 388,   37*2048+ 677,   10*2048+1055,    0*2048+1179,
   0*2048+ 278,   20*2048+ 516,    9*2048+ 952,    0*2048+1180,
   4*2048+  37,    0*2048+ 308,    9*2048+ 467,    0*2048+1181,
   0*2048+ 333,    5*2048+ 334,   33*2048+ 362,    0*2048+1182,
   8*2048+ 232,   24*2048+ 279,    0*2048+ 363,    0*2048+1183,
  26*2048+ 258,    0*2048+ 389,   36*2048+ 572,    0*2048+1184,
   0*2048+ 280,   43*2048+ 335,   27*2048+ 760,    0*2048+1185,
   0*2048+ 309,   25*2048+ 678,   35*2048+1030,    0*2048+1186,
   0*2048+ 336,   39*2048+ 390,   31*2048+ 843,    0*2048+1187,
  30*2048+  15,    0*2048+ 364,   13*2048+ 922,    0*2048+1188,
  37*2048+  66,    0*2048+ 391,   31*2048+ 439,    0*2048+1189,
  16*2048+  16,    0*2048+ 281,   12*2048+1031,    0*2048+1190,
   0*2048+ 310,   10*2048+ 844,   42*2048+ 923,    0*2048+1191,
   0*2048+ 337,    7*2048+ 392,   22*2048+ 761,    0*2048+1192,
  10*2048+  67,    0*2048+ 365,   14*2048+ 735,    0*2048+1193,
  29*2048+ 150,   14*2048+ 176,    0*2048+ 393,    0*2048+1194,
  16*2048+  38,    0*2048+ 282,   25*2048+ 283,    0*2048+1195,
   0*2048+ 311,   34*2048+ 492,   18*2048+ 601,    0*2048+1196,
   0*2048+ 338,   33*2048+ 493,    8*2048+ 517,    0*2048+1197,
  38*2048+ 151,    0*2048+ 366,   12*2048+ 976,    0*2048+1198,
   0*2048+ 394,   29*2048+ 602,   27*2048+ 924,    0*2048+1199,
   0*2048+ 412,   23*2048+ 575,   39*2048+ 895,    0*2048+1205,
   0*2048+ 441,   34*2048+ 790,   19*2048+ 870,    0*2048+1206,
   4*2048+ 177,    0*2048+ 470,   15*2048+ 625,    0*2048+1207,
  30*2048+ 284,    0*2048+ 496,    5*2048+ 680,    0*2048+1208,
   0*2048+ 519,   37*2048+ 520,   17*2048+ 736,    0*2048+1209,
  11*2048+  68,    0*2048+ 413,   12*2048+ 626,    0*2048+1210,
  21*2048+  95,    0*2048+ 442,   28*2048+ 521,    0*2048+1211,
  22*2048+ 259,    0*2048+ 471,   34*2048+ 576,    0*2048+1212,
  21*2048+ 285,    0*2048+ 497,   37*2048+ 953,    0*2048+1213,
   0*2048+ 522,   37*2048+ 845,   12*2048+1003,    0*2048+1214,
   0*2048+ 414,   25*2048+ 577,   42*2048+ 978,    0*2048+1215,
  29*2048+ 286,    0*2048+ 443,    2*2048+ 871,    0*2048+1216,
   0*2048+ 472,   35*2048+ 498,   16*2048+ 872,    0*2048+1217,
   0*2048+ 499,   36*2048+ 762,   15*2048+1057,    0*2048+1218,
  11*2048+ 122,    0*2048+ 523,   37*2048+ 814,    0*2048+1219,
  10*2048+  17,    0*2048+ 415,   20*2048+ 656,    0*2048+1220,
   4*2048+ 178,    0*2048+ 444,    9*2048+ 603,    0*2048+1221,
   0*2048+ 473,    5*2048+ 474,   33*2048+ 500,    0*2048+1222,
   8*2048+ 368,   24*2048+ 416,    0*2048+ 501,    0*2048+1223,
  26*2048+ 395,    0*2048+ 524,   36*2048+ 708,    0*2048+1224,
   0*2048+ 417,   43*2048+ 475,   27*2048+ 896,    0*2048+1225,
  36*2048+  96,    0*2048+ 445,   25*2048+ 815,    0*2048+1226,
   0*2048+ 476,   39*2048+ 525,   31*2048+ 979,    0*2048+1227,
  30*2048+ 152,    0*2048+ 502,   13*2048+1058,    0*2048+1228,
  37*2048+ 202,    0*2048+ 526,   31*2048+ 578,    0*2048+1229,
  13*2048+  97,   16*2048+ 153,    0*2048+ 418,    0*2048+1230,
   0*2048+ 446,   10*2048+ 980,   42*2048+1059,    0*2048+1231,
   0*2048+ 477,    7*2048+ 527,   22*2048+ 897,    0*2048+1232,
  10*2048+ 203,    0*2048+ 503,   14*2048+ 873,    0*2048+1233,
  29*2048+ 287,   14*2048+ 312,    0*2048+ 528,    0*2048+1234,
  16*2048+ 179,    0*2048+ 419,   25*2048+ 420,    0*2048+1235,
   0*2048+ 447,   34*2048+ 627,   18*2048+ 737,    0*2048+1236,
   0*2048+ 478,   33*2048+ 628,    8*2048+ 657,    0*2048+1237,
  13*2048+  39,   38*2048+ 288,    0*2048+ 504,    0*2048+1238,
   0*2048+ 529,   29*2048+ 738,   27*2048+1060,    0*2048+1239,
   0*2048+ 548,   23*2048+ 711,   39*2048+1032,    0*2048+1245,
   0*2048+ 580,   34*2048+ 926,   19*2048+1005,    0*2048+1246,
   4*2048+ 313,    0*2048+ 606,   15*2048+ 763,    0*2048+1247,
  30*2048+ 421,    0*2048+ 631,    5*2048+ 817,    0*2048+1248,
   0*2048+ 659,   37*2048+ 660,   17*2048+ 874,    0*2048+1249,
  11*2048+ 204,    0*2048+ 549,   12*2048+ 764,    0*2048+1250,
  21*2048+ 234,    0*2048+ 581,   28*2048+ 661,    0*2048+1251,
  22*2048+ 396,    0*2048+ 607,   34*2048+ 712,    0*2048+1252,
  38*2048+  18,   21*2048+ 422,    0*2048+ 632,    0*2048+1253,
  13*2048+  69,    0*2048+ 662,   37*2048+ 981,    0*2048+1254,
  43*2048+  41,    0*2048+ 550,   25*2048+ 713,    0*2048+1255,
  29*2048+ 423,    0*2048+ 582,    2*2048+1006,    0*2048+1256,
   0*2048+ 608,   35*2048+ 633,   16*2048+1007,    0*2048+1257,
  16*2048+ 124,    0*2048+ 634,   36*2048+ 898,    0*2048+1258,
  11*2048+ 260,    0*2048+ 663,   37*2048+ 954,    0*2048+1259,
  10*2048+ 154,    0*2048+ 551,   20*2048+ 792,    0*2048+1260,
   4*2048+ 314,    0*2048+ 583,    9*2048+ 739,    0*2048+1261,
   0*2048+ 609,    5*2048+ 610,   33*2048+ 635,    0*2048+1262,
   8*2048+ 506,   24*2048+ 552,    0*2048+ 636,    0*2048+1263,
  26*2048+ 530,    0*2048+ 664,   36*2048+ 846,    0*2048+1264,
   0*2048+ 553,   43*2048+ 611,   27*2048+1033,    0*2048+1265,
  36*2048+ 235,    0*2048+ 584,   25*2048+ 955,    0*2048+1266,
  32*2048+  42,    0*2048+ 612,   39*2048+ 665,    0*2048+1267,
  14*2048+ 125,   30*2048+ 289,    0*2048+ 637,    0*2048+1268,
  37*2048+ 340,    0*2048+ 666,   31*2048+ 714,    0*2048+1269,
  13*2048+ 236,   16*2048+ 290,    0*2048+ 554,    0*2048+1270,
  11*2048+  43,   43*2048+ 126,    0*2048+ 585,    0*2048+1271,
   0*2048+ 613,    7*2048+ 667,   22*2048+1034,    0*2048+1272,
  10*2048+ 341,    0*2048+ 638,   14*2048+1008,    0*2048+1273,
  29*2048+ 424,   14*2048+ 448,    0*2048+ 668,    0*2048+1274,
  16*2048+ 315,    0*2048+ 555,   25*2048+ 556,    0*2048+1275,
   0*2048+ 586,   34*2048+ 765,   18*2048+ 875,    0*2048+1276,
   0*2048+ 614,   33*2048+ 766,    8*2048+ 793,    0*2048+1277,
  13*2048+ 180,   38*2048+ 425,    0*2048+ 639,    0*2048+1278,
  28*2048+ 127,    0*2048+ 669,   29*2048+ 876,    0*2048+1279,
  40*2048+  98,    0*2048+ 684,   23*2048+ 849,    0*2048+1285,
  20*2048+  71,    0*2048+ 716,   34*2048+1062,    0*2048+1286,
   4*2048+ 449,    0*2048+ 742,   15*2048+ 899,    0*2048+1287,
  30*2048+ 557,    0*2048+ 769,    5*2048+ 957,    0*2048+1288,
   0*2048+ 795,   37*2048+ 796,   17*2048+1009,    0*2048+1289,
  11*2048+ 342,    0*2048+ 685,   12*2048+ 900,    0*2048+1290,
  21*2048+ 370,    0*2048+ 717,   28*2048+ 797,    0*2048+1291,
  22*2048+ 531,    0*2048+ 743,   34*2048+ 850,    0*2048+1292,
  38*2048+ 155,   21*2048+ 558,    0*2048+ 770,    0*2048+1293,
  38*2048+  44,   13*2048+ 205,    0*2048+ 798,    0*2048+1294,
  43*2048+ 182,    0*2048+ 686,   25*2048+ 851,    0*2048+1295,
   3*2048+  72,   29*2048+ 559,    0*2048+ 718,    0*2048+1296,
  17*2048+  73,    0*2048+ 744,   35*2048+ 771,    0*2048+1297,
  16*2048+ 262,    0*2048+ 772,   36*2048+1035,    0*2048+1298,
  38*2048+  19,   11*2048+ 397,    0*2048+ 799,    0*2048+1299,
  10*2048+ 291,    0*2048+ 687,   20*2048+ 928,    0*2048+1300,
   4*2048+ 450,    0*2048+ 719,    9*2048+ 877,    0*2048+1301,
   0*2048+ 745,    5*2048+ 746,   33*2048+ 773,    0*2048+1302,
   8*2048+ 641,   24*2048+ 688,    0*2048+ 774,    0*2048+1303,
  26*2048+ 670,    0*2048+ 800,   36*2048+ 982,    0*2048+1304,
  28*2048+  99,    0*2048+ 689,   43*2048+ 747,    0*2048+1305,
  26*2048+  20,   36*2048+ 371,    0*2048+ 720,    0*2048+1306,
  32*2048+ 183,    0*2048+ 748,   39*2048+ 801,    0*2048+1307,
  14*2048+ 263,   30*2048+ 426,    0*2048+ 775,    0*2048+1308,
  37*2048+ 480,    0*2048+ 802,   31*2048+ 852,    0*2048+1309,
  13*2048+ 372,   16*2048+ 427,    0*2048+ 690,    0*2048+1310,
  11*2048+ 184,   43*2048+ 264,    0*2048+ 721,    0*2048+1311,
  23*2048+ 100,    0*2048+ 749,    7*2048+ 803,    0*2048+1312,
  15*2048+  74,   10*2048+ 481,    0*2048+ 776,    0*2048+1313,
  29*2048+ 560,   14*2048+ 587,    0*2048+ 804,    0*2048+1314,
  16*2048+ 451,    0*2048+ 691,   25*2048+ 692,    0*2048+1315,
   0*2048+ 722,   34*2048+ 901,   18*2048+1010,    0*2048+1316,
   0*2048+ 750,   33*2048+ 902,    8*2048+ 929,    0*2048+1317,
  13*2048+ 316,   38*2048+ 561,    0*2048+ 777,    0*2048+1318,
  28*2048+ 265,    0*2048+ 805,   29*2048+1011,    0*2048+1319,
  40*2048+ 237,    0*2048+ 821,   23*2048+ 985,    0*2048+1325,
  35*2048+ 129,   20*2048+ 207,    0*2048+ 854,    0*2048+1326,
   4*2048+ 588,    0*2048+ 880,   15*2048+1036,    0*2048+1327,
   6*2048+  22,   30*2048+ 693,    0*2048+ 905,    0*2048+1328,
  18*2048+  75,    0*2048+ 931,   37*2048+ 932,    0*2048+1329,
  11*2048+ 482,    0*2048+ 822,   12*2048+1037,    0*2048+1330,
  21*2048+ 508,    0*2048+ 855,   28*2048+ 933,    0*2048+1331,
  22*2048+ 671,    0*2048+ 881,   34*2048+ 986,    0*2048+1332,
  38*2048+ 292,   21*2048+ 694,    0*2048+ 906,    0*2048+1333,
  38*2048+ 185,   13*2048+ 343,    0*2048+ 934,    0*2048+1334,
  43*2048+ 318,    0*2048+ 823,   25*2048+ 987,    0*2048+1335,
   3*2048+ 208,   29*2048+ 695,    0*2048+ 856,    0*2048+1336,
  17*2048+ 209,    0*2048+ 882,   35*2048+ 907,    0*2048+1337,
  37*2048+ 101,   16*2048+ 399,    0*2048+ 908,    0*2048+1338,
  38*2048+ 156,   11*2048+ 532,    0*2048+ 935,    0*2048+1339,
  10*2048+ 428,    0*2048+ 824,   20*2048+1064,    0*2048+1340,
   4*2048+ 589,    0*2048+ 857,    9*2048+1012,    0*2048+1341,
   0*2048+ 883,    5*2048+ 884,   33*2048+ 909,    0*2048+1342,
   8*2048+ 779,   24*2048+ 825,    0*2048+ 910,    0*2048+1343,
  37*2048+  45,   26*2048+ 806,    0*2048+ 936,    0*2048+1344,
  28*2048+ 238,    0*2048+ 826,   43*2048+ 885,    0*2048+1345,
  26*2048+ 157,   36*2048+ 509,    0*2048+ 858,    0*2048+1346,
  32*2048+ 319,    0*2048+ 886,   39*2048+ 937,    0*2048+1347,
  14*2048+ 400,   30*2048+ 562,    0*2048+ 911,    0*2048+1348,
  37*2048+ 616,    0*2048+ 938,   31*2048+ 988,    0*2048+1349,
  13*2048+ 510,   16*2048+ 563,    0*2048+ 827,    0*2048+1350,
  11*2048+ 320,   43*2048+ 401,    0*2048+ 859,    0*2048+1351,
  23*2048+ 239,    0*2048+ 887,    7*2048+ 939,    0*2048+1352,
  15*2048+ 210,   10*2048+ 617,    0*2048+ 912,    0*2048+1353,
  29*2048+ 696,   14*2048+ 723,    0*2048+ 940,    0*2048+1354,
  16*2048+ 590,    0*2048+ 828,   25*2048+ 829,    0*2048+1355,
  19*2048+  76,    0*2048+ 860,   34*2048+1038,    0*2048+1356,
   0*2048+ 888,   33*2048+1039,    8*2048+1065,    0*2048+1357,
  13*2048+ 452,   38*2048+ 697,    0*2048+ 913,    0*2048+1358,
  30*2048+  77,   28*2048+ 402,    0*2048+ 941,    0*2048+1359,
  24*2048+  48,   40*2048+ 373,    0*2048+ 961,    0*2048+1365,
  35*2048+ 267,   20*2048+ 345,    0*2048+ 990,    0*2048+1366,
  16*2048+ 102,    4*2048+ 724,    0*2048+1015,    0*2048+1367,
   6*2048+ 159,   30*2048+ 830,    0*2048+1042,    0*2048+1368,
  18*2048+ 211,    0*2048+1067,   37*2048+1068,    0*2048+1369,
  13*2048+ 103,   11*2048+ 618,    0*2048+ 962,    0*2048+1370,
  21*2048+ 643,    0*2048+ 991,   28*2048+1069,    0*2048+1371,
  35*2048+  49,   22*2048+ 807,    0*2048+1016,    0*2048+1372,
  38*2048+ 429,   21*2048+ 831,    0*2048+1043,    0*2048+1373,
  38*2048+ 321,   13*2048+ 483,    0*2048+1070,    0*2048+1374,
  26*2048+  50,   43*2048+ 454,    0*2048+ 963,    0*2048+1375,
   3*2048+ 346,   29*2048+ 832,    0*2048+ 992,    0*2048+1376,
  17*2048+ 347,    0*2048+1017,   35*2048+1044,    0*2048+1377,
  37*2048+ 240,   16*2048+ 534,    0*2048+1045,    0*2048+1378,
  38*2048+ 293,   11*2048+ 672,    0*2048+1071,    0*2048+1379,
  21*2048+ 131,   10*2048+ 564,    0*2048+ 964,    0*2048+1380,
  10*2048+  78,    4*2048+ 725,    0*2048+ 993,    0*2048+1381,
   0*2048+1018,    5*2048+1019,   33*2048+1046,    0*2048+1382,
   8*2048+ 915,   24*2048+ 965,    0*2048+1047,    0*2048+1383,
  37*2048+ 186,   26*2048+ 942,    0*2048+1072,    0*2048+1384,
  28*2048+ 374,    0*2048+ 966,   43*2048+1020,    0*2048+1385,
  26*2048+ 294,   36*2048+ 644,    0*2048+ 994,    0*2048+1386,
  32*2048+ 455,    0*2048+1021,   39*2048+1073,    0*2048+1387,
  14*2048+ 535,   30*2048+ 698,    0*2048+1048,    0*2048+1388,
  32*2048+  51,   37*2048+ 752,    0*2048+1074,    0*2048+1389,
  13*2048+ 645,   16*2048+ 699,    0*2048+ 967,    0*2048+1390,
  11*2048+ 456,   43*2048+ 536,    0*2048+ 995,    0*2048+1391,
  23*2048+ 375,    0*2048+1022,    7*2048+1075,    0*2048+1392,
  15*2048+ 348,   10*2048+ 753,    0*2048+1049,    0*2048+1393,
  29*2048+ 833,   14*2048+ 861,    0*2048+1076,    0*2048+1394,
  16*2048+ 726,    0*2048+ 968,   25*2048+ 969,    0*2048+1395,
  35*2048+ 104,   19*2048+ 212,    0*2048+ 996,    0*2048+1396,
  34*2048+ 105,    9*2048+ 132,    0*2048+1023,    0*2048+1397,
  13*2048+ 591,   38*2048+ 834,    0*2048+1050,    0*2048+1398,
  30*2048+ 213,   28*2048+ 537,    0*2048+1077,    0*2048+1399,
   0*2048+   0,   20*2048+ 135,   17*2048+ 864,   38*2048+1026,    0*2048+1080,
   0*2048+  27,   36*2048+ 270,   33*2048+ 459,   21*2048+ 891,    0*2048+1081,
   0*2048+  54,   28*2048+ 243,   43*2048+ 567,   29*2048+ 648,    0*2048+1082,
   0*2048+  81,   20*2048+ 162,   39*2048+ 163,    7*2048+ 378,    0*2048+1083,
  12*2048+  55,   23*2048+  82,    0*2048+ 108,   15*2048+ 136,    0*2048+1084,
  39*2048+  92,    0*2048+ 137,   20*2048+ 272,   17*2048+ 999,    0*2048+1120,
   0*2048+ 168,   36*2048+ 407,   33*2048+ 595,   21*2048+1028,    0*2048+1121,
   0*2048+ 190,   28*2048+ 380,   43*2048+ 703,   29*2048+ 784,    0*2048+1122,
   0*2048+ 220,   20*2048+ 298,   39*2048+ 299,    7*2048+ 513,    0*2048+1123,
  12*2048+ 191,   23*2048+ 221,    0*2048+ 246,   15*2048+ 273,    0*2048+1124,
  18*2048+  65,   39*2048+ 231,    0*2048+ 274,   20*2048+ 409,    0*2048+1160,
  22*2048+  94,    0*2048+ 304,   36*2048+ 543,   33*2048+ 731,    0*2048+1161,
   0*2048+ 328,   28*2048+ 515,   43*2048+ 841,   29*2048+ 920,    0*2048+1162,
   0*2048+ 356,   20*2048+ 434,   39*2048+ 435,    7*2048+ 653,    0*2048+1163,
  12*2048+ 329,   23*2048+ 357,    0*2048+ 383,   15*2048+ 410,    0*2048+1164,
  18*2048+ 201,   39*2048+ 367,    0*2048+ 411,   20*2048+ 545,    0*2048+1200,
  22*2048+ 233,    0*2048+ 440,   36*2048+ 679,   33*2048+ 869,    0*2048+1201,
   0*2048+ 468,   28*2048+ 655,   43*2048+ 977,   29*2048+1056,    0*2048+1202,
   0*2048+ 494,   20*2048+ 573,   39*2048+ 574,    7*2048+ 789,    0*2048+1203,
  12*2048+ 469,   23*2048+ 495,    0*2048+ 518,   15*2048+ 546,    0*2048+1204,
  18*2048+ 339,   39*2048+ 505,    0*2048+ 547,   20*2048+ 681,    0*2048+1240,
  22*2048+ 369,    0*2048+ 579,   36*2048+ 816,   33*2048+1004,    0*2048+1241,
  44*2048+  40,   30*2048+ 123,    0*2048+ 604,   28*2048+ 791,    0*2048+1242,
   0*2048+ 629,   20*2048+ 709,   39*2048+ 710,    7*2048+ 925,    0*2048+1243,
  12*2048+ 605,   23*2048+ 630,    0*2048+ 658,   15*2048+ 682,    0*2048+1244,
  18*2048+ 479,   39*2048+ 640,    0*2048+ 683,   20*2048+ 818,    0*2048+1280,
  34*2048+  70,   22*2048+ 507,    0*2048+ 715,   36*2048+ 956,    0*2048+1281,
  44*2048+ 181,   30*2048+ 261,    0*2048+ 740,   28*2048+ 927,    0*2048+1282,
   0*2048+ 767,   20*2048+ 847,   39*2048+ 848,    7*2048+1061,    0*2048+1283,
  12*2048+ 741,   23*2048+ 768,    0*2048+ 794,   15*2048+ 819,    0*2048+1284,
  18*2048+ 615,   39*2048+ 778,    0*2048+ 820,   20*2048+ 958,    0*2048+1320,
  37*2048+  21,   34*2048+ 206,   22*2048+ 642,    0*2048+ 853,    0*2048+1321,
  44*2048+ 317,   30*2048+ 398,    0*2048+ 878,   28*2048+1063,    0*2048+1322,
   8*2048+ 128,    0*2048+ 903,   20*2048+ 983,   39*2048+ 984,    0*2048+1323,
  12*2048+ 879,   23*2048+ 904,    0*2048+ 930,   15*2048+ 959,    0*2048+1324,
  21*2048+  23,   18*2048+ 751,   39*2048+ 914,    0*2048+ 960,    0*2048+1360,
  37*2048+ 158,   34*2048+ 344,   22*2048+ 780,    0*2048+ 989,    0*2048+1361,
  29*2048+ 130,   44*2048+ 453,   30*2048+ 533,    0*2048+1013,    0*2048+1362,
  21*2048+  46,   40*2048+  47,    8*2048+ 266,    0*2048+1040,    0*2048+1363,
  16*2048+  24,   12*2048+1014,   23*2048+1041,    0*2048+1066,    0*2048+1364);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if RdAddr < ROM'length then
				Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , Do'length );
			end if;
		end if;
	end process;

end Behavioral;