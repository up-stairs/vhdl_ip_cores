LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VNP_Input_Edge_Memory is
	Port (
		clk			: in  std_logic;
		
		RdAddr		: in  std_logic_vector(13 downto 0);
		Do			: out std_logic_vector(11 downto 0)
	);
end VNP_Input_Edge_Memory;

architecture Behavioral of VNP_Input_Edge_Memory is	
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 15272-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
   2,    6, 2048+1152,
   7,   10, 2048+1153,
  11,   14, 2048+1154,
  15,   18, 2048+1155,
  19,   22, 2048+1156,
  23,   25, 2048+1157,
  26,   29, 2048+1158,
  30,   33, 2048+1159,
  34,   37, 2048+1160,
  38,   41, 2048+1161,
  42,   45, 2048+1162,
  46,   49, 2048+1163,
  50,   52, 2048+1164,
  53,   55, 2048+1165,
  56,   58, 2048+1166,
  59,   62, 2048+1167,
  63,   66, 2048+1168,
  67,   70, 2048+1169,
  71,   74, 2048+1170,
  75,   77, 2048+1171,
  78,   81, 2048+1172,
  82,   85, 2048+1173,
  86,   89, 2048+1174,
  90,   93, 2048+1175,
  94,   97, 2048+1176,
  98,  100, 2048+1177,
 101,  103, 2048+1178,
 104,  106, 2048+1179,
 107,  110, 2048+1180,
 111,  113, 2048+1181,
 114,  117, 2048+1182,
 118,  121, 2048+1183,
 122,  125, 2048+1184,
 126,  129, 2048+1185,
 130,  133, 2048+1186,
 134,  137, 2048+1187,
 138,  141, 2048+1188,
 142,  145, 2048+1189,
 146,  149, 2048+1190,
 150,  153, 2048+1191,
 154,  157, 2048+1192,
 158,  160, 2048+1193,
 161,  164, 2048+1194,
 165,  168, 2048+1195,
 169,  172, 2048+1196,
 173,  176, 2048+1197,
 177,  180, 2048+1198,
 181,  184, 2048+1199,
 185,  187, 2048+1200,
 188,  190, 2048+1201,
 191,  193, 2048+1202,
 194,  197, 2048+1203,
 198,  201, 2048+1204,
 202,  205, 2048+1205,
 206,  209, 2048+1206,
 210,  212, 2048+1207,
 213,  216, 2048+1208,
 217,  220, 2048+1209,
 221,  224, 2048+1210,
 225,  228, 2048+1211,
 229,  232, 2048+1212,
 233,  235, 2048+1213,
 236,  238, 2048+1214,
 239,  241, 2048+1215,
 242,  245, 2048+1216,
 246,  248, 2048+1217,
 249,  252, 2048+1218,
 253,  256, 2048+1219,
 257,  260, 2048+1220,
 261,  264, 2048+1221,
 265,  268, 2048+1222,
 269,  272, 2048+1223,
 273,  276, 2048+1224,
 277,  280, 2048+1225,
 281,  284, 2048+1226,
 285,  288, 2048+1227,
 289,  292, 2048+1228,
 293,  295, 2048+1229,
 296,  299, 2048+1230,
 300,  303, 2048+1231,
 304,  307, 2048+1232,
 308,  311, 2048+1233,
 312,  315, 2048+1234,
 316,  319, 2048+1235,
 320,  322, 2048+1236,
 323,  325, 2048+1237,
 326,  328, 2048+1238,
 329,  332, 2048+1239,
 333,  336, 2048+1240,
 337,  340, 2048+1241,
 341,  344, 2048+1242,
 345,  347, 2048+1243,
 348,  351, 2048+1244,
 352,  355, 2048+1245,
 356,  359, 2048+1246,
 360,  363, 2048+1247,
 364,  367, 2048+1248,
 368,  370, 2048+1249,
 371,  373, 2048+1250,
 374,  376, 2048+1251,
 377,  380, 2048+1252,
 381,  383, 2048+1253,
 384,  387, 2048+1254,
 388,  391, 2048+1255,
 392,  395, 2048+1256,
 396,  399, 2048+1257,
 400,  403, 2048+1258,
 404,  407, 2048+1259,
 408,  411, 2048+1260,
 412,  415, 2048+1261,
 416,  419, 2048+1262,
 420,  423, 2048+1263,
 424,  427, 2048+1264,
 428,  430, 2048+1265,
 431,  434, 2048+1266,
 435,  438, 2048+1267,
 439,  442, 2048+1268,
 443,  446, 2048+1269,
 447,  450, 2048+1270,
 451,  454, 2048+1271,
 455,  457, 2048+1272,
 458,  460, 2048+1273,
 461,  463, 2048+1274,
 464,  467, 2048+1275,
 468,  471, 2048+1276,
 472,  475, 2048+1277,
 476,  479, 2048+1278,
 480,  482, 2048+1279,
 483,  486, 2048+1280,
 487,  490, 2048+1281,
 491,  494, 2048+1282,
 495,  498, 2048+1283,
 499,  502, 2048+1284,
 503,  505, 2048+1285,
 506,  508, 2048+1286,
 509,  511, 2048+1287,
 512,  515, 2048+1288,
 516,  518, 2048+1289,
 519,  522, 2048+1290,
 523,  526, 2048+1291,
 527,  530, 2048+1292,
 531,  534, 2048+1293,
 535,  538, 2048+1294,
 539,  542, 2048+1295,
 543,  546, 2048+1296,
 547,  550, 2048+1297,
 551,  554, 2048+1298,
 555,  558, 2048+1299,
 559,  562, 2048+1300,
 563,  565, 2048+1301,
 566,  569, 2048+1302,
 570,  573, 2048+1303,
 574,  577, 2048+1304,
 578,  581, 2048+1305,
 582,  585, 2048+1306,
 586,  589, 2048+1307,
 590,  592, 2048+1308,
 593,  595, 2048+1309,
 596,  598, 2048+1310,
 599,  602, 2048+1311,
 603,  606, 2048+1312,
 607,  610, 2048+1313,
 611,  614, 2048+1314,
 615,  617, 2048+1315,
 618,  621, 2048+1316,
 622,  625, 2048+1317,
 626,  629, 2048+1318,
 630,  633, 2048+1319,
 634,  637, 2048+1320,
 638,  640, 2048+1321,
 641,  643, 2048+1322,
 644,  646, 2048+1323,
 647,  650, 2048+1324,
 651,  653, 2048+1325,
 654,  657, 2048+1326,
 658,  661, 2048+1327,
 662,  665, 2048+1328,
 666,  669, 2048+1329,
 670,  673, 2048+1330,
 674,  677, 2048+1331,
 678,  681, 2048+1332,
 682,  685, 2048+1333,
 686,  689, 2048+1334,
 690,  693, 2048+1335,
 694,  697, 2048+1336,
 698,  700, 2048+1337,
 701,  704, 2048+1338,
 705,  708, 2048+1339,
 709,  712, 2048+1340,
 713,  716, 2048+1341,
 717,  720, 2048+1342,
 721,  724, 2048+1343,
 725,  727, 2048+1344,
 728,  730, 2048+1345,
 731,  733, 2048+1346,
 734,  737, 2048+1347,
 738,  741, 2048+1348,
 742,  745, 2048+1349,
 746,  749, 2048+1350,
 750,  752, 2048+1351,
 753,  756, 2048+1352,
 757,  760, 2048+1353,
 761,  764, 2048+1354,
 765,  768, 2048+1355,
 769,  772, 2048+1356,
 773,  775, 2048+1357,
 776,  778, 2048+1358,
 779,  781, 2048+1359,
 782,  785, 2048+1360,
 786,  788, 2048+1361,
 789,  792, 2048+1362,
 793,  796, 2048+1363,
 797,  800, 2048+1364,
 801,  804, 2048+1365,
 805,  808, 2048+1366,
 809,  812, 2048+1367,
 813,  816, 2048+1368,
 817,  820, 2048+1369,
 821,  824, 2048+1370,
 825,  828, 2048+1371,
 829,  832, 2048+1372,
 833,  835, 2048+1373,
 836,  839, 2048+1374,
 840,  843, 2048+1375,
 844,  847, 2048+1376,
 848,  851, 2048+1377,
 852,  855, 2048+1378,
 856,  859, 2048+1379,
 860,  862, 2048+1380,
 863,  865, 2048+1381,
 866,  868, 2048+1382,
 869,  872, 2048+1383,
 873,  876, 2048+1384,
 877,  880, 2048+1385,
 881,  884, 2048+1386,
 885,  887, 2048+1387,
 888,  891, 2048+1388,
 892,  895, 2048+1389,
 896,  899, 2048+1390,
 900,  903, 2048+1391,
 904,  907, 2048+1392,
 908,  910, 2048+1393,
 911,  913, 2048+1394,
 914,  916, 2048+1395,
 917,  920, 2048+1396,
 921,  923, 2048+1397,
 924,  927, 2048+1398,
 928,  931, 2048+1399,
 932,  935, 2048+1400,
 936,  939, 2048+1401,
 940,  943, 2048+1402,
 944,  947, 2048+1403,
 948,  951, 2048+1404,
 952,  955, 2048+1405,
 956,  959, 2048+1406,
 960,  963, 2048+1407,
 964,  967, 2048+1408,
 968,  970, 2048+1409,
 971,  974, 2048+1410,
 975,  978, 2048+1411,
 979,  982, 2048+1412,
 983,  986, 2048+1413,
 987,  990, 2048+1414,
 991,  994, 2048+1415,
 995,  997, 2048+1416,
 998, 1000, 2048+1417,
1001, 1003, 2048+1418,
1004, 1007, 2048+1419,
1008, 1011, 2048+1420,
1012, 1015, 2048+1421,
1016, 1019, 2048+1422,
1020, 1022, 2048+1423,
1023, 1026, 2048+1424,
1027, 1030, 2048+1425,
1031, 1034, 2048+1426,
1035, 1038, 2048+1427,
1039, 1042, 2048+1428,
1043, 1045, 2048+1429,
1046, 1048, 2048+1430,
1049, 1051, 2048+1431,
1052, 1055, 2048+1432,
1056, 1058, 2048+1433,
1059, 1062, 2048+1434,
1063, 1066, 2048+1435,
1067, 1070, 2048+1436,
1071, 1074, 2048+1437,
1075, 1078, 2048+1438,
   3, 1079, 2048+1439,
 254,  440,  748, 2048+1084,
 743,  814, 1032, 2048+1085,
 398,  758,  780, 2048+1086,
 148,  528,  783, 2048+1087,
 182,  203,  305, 2048+1088,
 389,  575,  883, 2048+1093,
  87,  878,  949, 2048+1094,
 533,  893,  915, 2048+1095,
 283,  663,  918, 2048+1096,
 317,  338,  441, 2048+1097,
 524,  710, 1018, 2048+1102,
   4,  222, 1013, 2048+1103,
 668, 1028, 1050, 2048+1104,
 418,  798, 1053, 2048+1105,
 452,  473,  576, 2048+1106,
  73,  660,  845, 2048+1111,
  68,  139,  358, 2048+1112,
  83,  105,  803, 2048+1113,
 108,  553,  933, 2048+1114,
 587,  608,  711, 2048+1115,
 208,  795,  980, 2048+1120,
 204,  274,  493, 2048+1121,
 218,  240,  938, 2048+1122,
 243,  688, 1068, 2048+1123,
 722,  744,  846, 2048+1124,
  35,  343,  930, 2048+1129,
 339,  409,  628, 2048+1130,
 353,  375, 1073, 2048+1131,
 123,  378,  823, 2048+1132,
 857,  879,  981, 2048+1133,
 170,  478, 1065, 2048+1138,
 474,  544,  763, 2048+1139,
 128,  488,  510, 2048+1140,
 259,  513,  958, 2048+1141,
  36,  992, 1014, 2048+1142,
 120,  306,  613, 2048+1147,
 609,  680,  898, 2048+1148,
 263,  624,  645, 2048+1149,
  13,  394,  649, 2048+1150,
  48,   69,  171, 2048+1151,
  43,   60,  151,  357,  459,  540,  648,  777,  826,  867,  925,  972, 2048+1080,
  20,  131,  143,  346,  432,  548,  718,  747,  766,  870,  874, 1044, 2048+1081,
  91,  147,  309,  349,  397,  444,  591,  635,  706,  875,  926,  976, 2048+1082,
  47,  132,  230,  258,  294,  350,  623,  659,  679,  830,  945, 1057, 2048+1083,
  27,  178,  195,  286,  492,  594,  675,  784,  912,  961, 1002, 1060, 2048+1089,
  99,  155,  266,  278,  481,  567,  683,  853,  882,  901, 1005, 1009, 2048+1090,
  31,  226,  282,  445,  484,  532,  579,  726,  770,  841, 1010, 1061, 2048+1091,
   0,  112,  183,  267,  365,  393,  429,  485,  759,  794,  815,  965, 2048+1092,
  16,   57,  115,  162,  313,  330,  421,  627,  729,  810,  919, 1047, 2048+1098,
  61,   64,  234,  290,  401,  413,  616,  702,  818,  988, 1017, 1036, 2048+1099,
  65,  116,  166,  361,  417,  580,  619,  667,  714,  861,  905,  977, 2048+1100,
  21,  135,  247,  318,  402,  500,  529,  564,  620,  894,  929,  950, 2048+1101,
 102,  152,  192,  250,  297,  448,  465,  556,  762,  864,  946, 1054, 2048+1107,
  44,   72,   92,  196,  199,  369,  425,  536,  549,  751,  837,  953, 2048+1108,
  32,  200,  251,  301,  496,  552,  715,  754,  802,  849,  996, 1040, 2048+1109,
   5,  156,  270,  382,  453,  537,  636,  664,  699,  755, 1029, 1064, 2048+1110,
   1,  109,  237,  287,  327,  385,  433,  583,  600,  691,  897,  999, 2048+1116,
   8,  179,  207,  227,  331,  334,  504,  560,  671,  684,  886,  973, 2048+1117,
  51,   95,  167,  335,  386,  436,  631,  687,  850,  889,  937,  984, 2048+1118,
  84,  119,  140,  291,  405,  517,  588,  672,  771,  799,  834,  890, 2048+1119,
  54,  136,  244,  372,  422,  462,  520,  568,  719,  735,  827, 1033, 2048+1125,
  28,  144,  314,  342,  362,  466,  469,  639,  695,  806,  819, 1021, 2048+1126,
  39,  186,  231,  302,  470,  521,  571,  767,  822,  985, 1024, 1072, 2048+1127,
 219,  255,  275,  426,  541,  652,  723,  807,  906,  934,  969, 1025, 2048+1128,
  88,  189,  271,  379,  507,  557,  597,  655,  703,  854,  871,  962, 2048+1134,
  76,  163,  279,  449,  477,  497,  601,  604,  774,  831,  941,  954, 2048+1135,
  40,   79,  127,  174,  321,  366,  437,  605,  656,  707,  902,  957, 2048+1136,
  24,   80,  354,  390,  410,  561,  676,  787,  858,  942, 1041, 1069, 2048+1137,
  17,  223,  324,  406,  514,  642,  692,  732,  790,  838,  989, 1006, 2048+1143,
   9,  211,  298,  414,  584,  612,  632,  736,  739,  909,  966, 1076, 2048+1144,
  12,  175,  214,  262,  310,  456,  501,  572,  740,  791,  842, 1037, 2048+1145,
  96,  124,  159,  215,  489,  525,  545,  696,  811,  922,  993, 1077, 2048+1146,

   3,    8, 2048+1320,
   9,   13, 2048+1321,
  14,   18, 2048+1322,
  19,   23, 2048+1323,
  24,   28, 2048+1324,
  29,   33, 2048+1325,
  34,   38, 2048+1326,
  39,   43, 2048+1327,
  44,   48, 2048+1328,
  49,   53, 2048+1329,
  54,   58, 2048+1330,
  59,   63, 2048+1331,
  64,   68, 2048+1332,
  69,   73, 2048+1333,
  74,   78, 2048+1334,
  79,   83, 2048+1335,
  84,   88, 2048+1336,
  89,   93, 2048+1337,
  94,   98, 2048+1338,
  99,  103, 2048+1339,
 104,  108, 2048+1340,
 109,  113, 2048+1341,
 114,  118, 2048+1342,
 119,  123, 2048+1343,
 124,  128, 2048+1344,
 129,  133, 2048+1345,
 134,  138, 2048+1346,
 139,  143, 2048+1347,
 144,  148, 2048+1348,
 149,  153, 2048+1349,
 154,  158, 2048+1350,
 159,  163, 2048+1351,
 164,  168, 2048+1352,
 169,  173, 2048+1353,
 174,  178, 2048+1354,
 179,  183, 2048+1355,
 184,  188, 2048+1356,
 189,  193, 2048+1357,
 194,  198, 2048+1358,
 199,  203, 2048+1359,
 204,  208, 2048+1360,
 209,  213, 2048+1361,
 214,  218, 2048+1362,
 219,  223, 2048+1363,
 224,  228, 2048+1364,
 229,  233, 2048+1365,
 234,  238, 2048+1366,
 239,  243, 2048+1367,
 244,  248, 2048+1368,
 249,  253, 2048+1369,
 254,  258, 2048+1370,
 259,  263, 2048+1371,
 264,  268, 2048+1372,
 269,  273, 2048+1373,
 274,  278, 2048+1374,
 279,  283, 2048+1375,
 284,  288, 2048+1376,
 289,  293, 2048+1377,
 294,  298, 2048+1378,
 299,  303, 2048+1379,
 304,  308, 2048+1380,
 309,  313, 2048+1381,
 314,  318, 2048+1382,
 319,  323, 2048+1383,
 324,  328, 2048+1384,
 329,  333, 2048+1385,
 334,  338, 2048+1386,
 339,  343, 2048+1387,
 344,  348, 2048+1388,
 349,  353, 2048+1389,
 354,  358, 2048+1390,
 359,  363, 2048+1391,
 364,  368, 2048+1392,
 369,  373, 2048+1393,
 374,  378, 2048+1394,
 379,  383, 2048+1395,
 384,  388, 2048+1396,
 389,  393, 2048+1397,
 394,  398, 2048+1398,
 399,  403, 2048+1399,
 404,  408, 2048+1400,
 409,  413, 2048+1401,
 414,  418, 2048+1402,
 419,  423, 2048+1403,
 424,  428, 2048+1404,
 429,  433, 2048+1405,
 434,  438, 2048+1406,
 439,  443, 2048+1407,
 444,  448, 2048+1408,
 449,  453, 2048+1409,
 454,  458, 2048+1410,
 459,  463, 2048+1411,
 464,  468, 2048+1412,
 469,  473, 2048+1413,
 474,  478, 2048+1414,
 479,  483, 2048+1415,
 484,  488, 2048+1416,
 489,  493, 2048+1417,
 494,  498, 2048+1418,
 499,  503, 2048+1419,
 504,  508, 2048+1420,
 509,  513, 2048+1421,
 514,  518, 2048+1422,
 519,  523, 2048+1423,
 524,  528, 2048+1424,
 529,  533, 2048+1425,
 534,  538, 2048+1426,
 539,  543, 2048+1427,
 544,  548, 2048+1428,
 549,  553, 2048+1429,
 554,  558, 2048+1430,
 559,  563, 2048+1431,
 564,  568, 2048+1432,
 569,  573, 2048+1433,
 574,  578, 2048+1434,
 579,  583, 2048+1435,
 584,  588, 2048+1436,
 589,  593, 2048+1437,
 594,  598, 2048+1438,
 599,  603, 2048+1439,
 604,  608, 2048+1440,
 609,  613, 2048+1441,
 614,  618, 2048+1442,
 619,  623, 2048+1443,
 624,  628, 2048+1444,
 629,  633, 2048+1445,
 634,  638, 2048+1446,
 639,  643, 2048+1447,
 644,  648, 2048+1448,
 649,  653, 2048+1449,
 654,  658, 2048+1450,
 659,  663, 2048+1451,
 664,  668, 2048+1452,
 669,  673, 2048+1453,
 674,  678, 2048+1454,
 679,  683, 2048+1455,
 684,  688, 2048+1456,
 689,  693, 2048+1457,
 694,  698, 2048+1458,
 699,  703, 2048+1459,
 704,  708, 2048+1460,
 709,  713, 2048+1461,
 714,  718, 2048+1462,
 719,  723, 2048+1463,
 724,  728, 2048+1464,
 729,  733, 2048+1465,
 734,  738, 2048+1466,
 739,  743, 2048+1467,
 744,  748, 2048+1468,
 749,  753, 2048+1469,
 754,  758, 2048+1470,
 759,  763, 2048+1471,
 764,  768, 2048+1472,
 769,  773, 2048+1473,
 774,  778, 2048+1474,
 779,  783, 2048+1475,
 784,  788, 2048+1476,
 789,  793, 2048+1477,
 794,  798, 2048+1478,
 799,  803, 2048+1479,
 804,  808, 2048+1480,
 809,  813, 2048+1481,
 814,  818, 2048+1482,
 819,  823, 2048+1483,
 824,  828, 2048+1484,
 829,  833, 2048+1485,
 834,  838, 2048+1486,
 839,  843, 2048+1487,
 844,  848, 2048+1488,
 849,  853, 2048+1489,
 854,  858, 2048+1490,
 859,  863, 2048+1491,
 864,  868, 2048+1492,
 869,  873, 2048+1493,
 874,  878, 2048+1494,
 879,  883, 2048+1495,
 884,  888, 2048+1496,
 889,  893, 2048+1497,
 894,  898, 2048+1498,
 899,  903, 2048+1499,
 904,  908, 2048+1500,
 909,  913, 2048+1501,
 914,  918, 2048+1502,
 919,  923, 2048+1503,
 924,  928, 2048+1504,
 929,  933, 2048+1505,
 934,  938, 2048+1506,
 939,  943, 2048+1507,
 944,  948, 2048+1508,
 949,  953, 2048+1509,
 954,  958, 2048+1510,
 959,  963, 2048+1511,
 964,  968, 2048+1512,
 969,  973, 2048+1513,
 974,  978, 2048+1514,
 979,  983, 2048+1515,
 984,  988, 2048+1516,
 989,  993, 2048+1517,
 994,  998, 2048+1518,
 999, 1003, 2048+1519,
1004, 1008, 2048+1520,
1009, 1013, 2048+1521,
1014, 1018, 2048+1522,
1019, 1023, 2048+1523,
1024, 1028, 2048+1524,
1029, 1033, 2048+1525,
1034, 1038, 2048+1526,
1039, 1043, 2048+1527,
1044, 1048, 2048+1528,
1049, 1053, 2048+1529,
1054, 1058, 2048+1530,
1059, 1063, 2048+1531,
1064, 1068, 2048+1532,
1069, 1073, 2048+1533,
1074, 1078, 2048+1534,
1079, 1083, 2048+1535,
1084, 1088, 2048+1536,
1089, 1093, 2048+1537,
1094, 1098, 2048+1538,
1099, 1103, 2048+1539,
1104, 1108, 2048+1540,
1109, 1113, 2048+1541,
1114, 1118, 2048+1542,
1119, 1123, 2048+1543,
1124, 1128, 2048+1544,
1129, 1133, 2048+1545,
1134, 1138, 2048+1546,
1139, 1143, 2048+1547,
1144, 1148, 2048+1548,
1149, 1153, 2048+1549,
1154, 1158, 2048+1550,
1159, 1163, 2048+1551,
1164, 1168, 2048+1552,
1169, 1173, 2048+1553,
1174, 1178, 2048+1554,
1179, 1183, 2048+1555,
1184, 1188, 2048+1556,
1189, 1193, 2048+1557,
1194, 1198, 2048+1558,
   4, 1199, 2048+1559,
 325,  491,  810, 2048+1205,
 551,  715, 1060, 2048+1206,
 406,  505,  725, 2048+1207,
 146,  950,  971, 2048+1208,
 111,  140,  615, 2048+1209,
  90,  450, 1170, 2048+1210,
  45,  220,  336, 2048+1211,
 170,  586,  815, 2048+1212,
 190,  885, 1040, 2048+1213,
 235,  535, 1070, 2048+1214,
 475,  641,  962, 2048+1220,
  10,  702,  865, 2048+1221,
 556,  657,  876, 2048+1222,
 296, 1100, 1121, 2048+1223,
 261,  290,  765, 2048+1224,
 121,  240,  600, 2048+1225,
 195,  370,  486, 2048+1226,
 320,  736,  966, 2048+1227,
 340, 1035, 1190, 2048+1228,
  20,  386,  685, 2048+1229,
 625,  791, 1112, 2048+1235,
 161,  852, 1015, 2048+1236,
 706,  807, 1027, 2048+1237,
  50,   71,  446, 2048+1238,
 411,  441,  915, 2048+1239,
 271,  390,  750, 2048+1240,
 345,  520,  636, 2048+1241,
 470,  887, 1116, 2048+1242,
 141,  492, 1185, 2048+1243,
 171,  537,  835, 2048+1244,
  62,  775,  941, 2048+1250,
 311, 1002, 1165, 2048+1251,
 856,  957, 1177, 2048+1252,
 200,  222,  596, 2048+1253,
 561,  591, 1065, 2048+1254,
 421,  540,  900, 2048+1255,
 496,  670,  787, 2048+1256,
  66,  620, 1037, 2048+1257,
 135,  291,  642, 2048+1258,
 321,  687,  985, 2048+1259,
 212,  925, 1091, 2048+1265,
 117,  461, 1152, 2048+1266,
 127, 1006, 1107, 2048+1267,
 350,  372,  746, 2048+1268,
  16,  711,  741, 2048+1269,
 571,  691, 1051, 2048+1270,
 646,  820,  937, 2048+1271,
 216,  771, 1187, 2048+1272,
 285,  442,  792, 2048+1273,
 471,  837, 1135, 2048+1274,
  41,  362, 1077, 2048+1280,
 102,  267,  611, 2048+1281,
  57,  277, 1156, 2048+1282,
 501,  522,  896, 2048+1283,
 166,  861,  891, 2048+1284,
   2,  721,  842, 2048+1285,
 796,  972, 1087, 2048+1286,
 137,  366,  921, 2048+1287,
 435,  592,  942, 2048+1288,
  85,  621,  987, 2048+1289,
  27,  192,  512, 2048+1295,
 252,  417,  762, 2048+1296,
 107,  207,  427, 2048+1297,
 651,  672, 1047, 2048+1298,
 316, 1011, 1042, 2048+1299,
 152,  871,  992, 2048+1300,
  37,  946, 1122, 2048+1301,
 287,  517, 1072, 2048+1302,
 587,  742, 1092, 2048+1303,
 236,  772, 1137, 2048+1304,
 177,  342,  662, 2048+1310,
 402,  567,  912, 2048+1311,
 257,  357,  577, 2048+1312,
 802,  822, 1197, 2048+1313,
 467, 1162, 1192, 2048+1314,
 302, 1022, 1142, 2048+1315,
  72,  187, 1097, 2048+1316,
  22,  437,  667, 2048+1317,
  42,  737,  892, 2048+1318,
  87,  387,  922, 2048+1319,
  15,  145,  160,  380,  480,  800,  825,  845,  880,  960,  965, 1160, 2048+1200,
  95,  155,  330,  385,  440,  490,  655,  690,  780,  961, 1025, 1075, 2048+1201,
 115,  120,  225,  335,  495,  656,  770,  840,  881,  970, 1050, 1095, 2048+1202,
   0,  105,  110,  116,  381,  465,  500,  585,  700,  785,  875, 1076, 2048+1203,
 375,  395,  405,  515,  550,  730,  755,  756,  760, 1020, 1045, 1130, 2048+1204,
 112,  165,  295,  310,  530,  630,  951,  975,  995, 1030, 1110, 1115, 2048+1215,
  25,  245,  305,  481,  536,  590,  640,  805,  841,  930, 1111, 1175, 2048+1216,
   1,   46,  265,  270,  376,  485,  645,  806,  920,  990, 1031, 1120, 2048+1217,
  26,  150,  255,  260,  266,  531,  616,  650,  735,  850,  935, 1026, 2048+1218,
  80,  525,  545,  555,  665,  701,  882,  905,  906,  910, 1171, 1195, 2048+1219,
  60,   65,  262,  315,  445,  460,  680,  781, 1101, 1125, 1145, 1180, 2048+1230,
  61,  125,  175,  396,  455,  631,  686,  740,  790,  955,  991, 1080, 2048+1231,
  70,  151,  196,  415,  420,  526,  635,  795,  956, 1071, 1140, 1181, 2048+1232,
 176,  300,  407,  410,  416,  681,  766,  801,  886, 1000, 1085, 1176, 2048+1233,
 122,  147,  230,  675,  695,  705,  816,  851, 1032, 1055, 1056, 1061, 2048+1234,
  51,   75,   96,  130,  210,  215,  412,  466,  595,  610,  830,  931, 2048+1245,
  30,  211,  275,  326,  546,  605,  782,  836,  890,  940, 1105, 1141, 2048+1246,
  21,   91,  131,  221,  301,  346,  565,  570,  676,  786,  945, 1106, 2048+1247,
  35,  126,  327,  451,  557,  560,  566,  831,  916,  952, 1036, 1150, 2048+1248,
   5,    6,   11,  272,  297,  382,  826,  846,  855,  967, 1001, 1182, 2048+1249,
 201,  226,  246,  280,  360,  365,  562,  617,  745,  761,  980, 1081, 2048+1260,
  55,   92,  180,  361,  425,  476,  696,  757,  932,  986, 1041, 1090, 2048+1261,
  56,  172,  241,  281,  371,  452,  497,  716,  720,  827,  936, 1096, 2048+1262,
 100,  185,  276,  477,  601,  707,  710,  717,  981, 1066, 1102, 1186, 2048+1263,
 132,  156,  157,  162,  422,  447,  532,  976,  996, 1005, 1117, 1151, 2048+1264,
  31,  351,  377,  397,  430,  510,  516,  712,  767,  895,  911, 1131, 2048+1275,
  40,  205,  242,  331,  511,  575,  626,  847,  907, 1082, 1136, 1191, 2048+1276,
  47,  206,  322,  391,  431,  521,  602,  647,  866,  870,  977, 1086, 2048+1277,
  17,   52,  136,  250,  337,  426,  627,  751,  857,  860,  867, 1132, 2048+1278,
  67,  101,  282,  306,  307,  312,  572,  597,  682, 1126, 1146, 1155, 2048+1279,
  81,  181,  502,  527,  547,  580,  660,  666,  862,  917, 1046, 1062, 2048+1290,
  32,   86,  142,  191,  355,  392,  482,  661,  726,  776,  997, 1057, 2048+1291,
  36,  197,  356,  472,  541,  581,  671,  752,  797, 1016, 1021, 1127, 2048+1292,
  82,  167,  202,  286,  400,  487,  576,  777,  901, 1007, 1010, 1017, 2048+1293,
  76,   97,  106,  217,  251,  432,  456,  457,  462,  722,  747,  832, 2048+1294,
  12,  231,  332,  652,  677,  697,  731,  811,  817, 1012, 1067, 1196, 2048+1305,
   7,  182,  237,  292,  341,  506,  542,  632,  812,  877,  926, 1147, 2048+1306,
  77,  186,  347,  507,  622,  692,  732,  821,  902,  947, 1166, 1172, 2048+1307,
 232,  317,  352,  436,  552,  637,  727,  927, 1052, 1157, 1161, 1167, 2048+1308,
 227,  247,  256,  367,  401,  582,  606,  607,  612,  872,  897,  982, 2048+1309,

   4,   10, 2048+1440,
  11,   16, 2048+1441,
  17,   22, 2048+1442,
  23,   28, 2048+1443,
  29,   34, 2048+1444,
  35,   40, 2048+1445,
  41,   46, 2048+1446,
  47,   52, 2048+1447,
  53,   58, 2048+1448,
  59,   64, 2048+1449,
  65,   70, 2048+1450,
  71,   76, 2048+1451,
  77,   82, 2048+1452,
  83,   88, 2048+1453,
  89,   94, 2048+1454,
  95,  100, 2048+1455,
 101,  106, 2048+1456,
 107,  112, 2048+1457,
 113,  118, 2048+1458,
 119,  124, 2048+1459,
 125,  130, 2048+1460,
 131,  136, 2048+1461,
 137,  142, 2048+1462,
 143,  148, 2048+1463,
 149,  154, 2048+1464,
 155,  160, 2048+1465,
 161,  166, 2048+1466,
 167,  172, 2048+1467,
 173,  178, 2048+1468,
 179,  184, 2048+1469,
 185,  190, 2048+1470,
 191,  196, 2048+1471,
 197,  202, 2048+1472,
 203,  208, 2048+1473,
 209,  214, 2048+1474,
 215,  220, 2048+1475,
 221,  226, 2048+1476,
 227,  232, 2048+1477,
 233,  238, 2048+1478,
 239,  244, 2048+1479,
 245,  250, 2048+1480,
 251,  256, 2048+1481,
 257,  262, 2048+1482,
 263,  268, 2048+1483,
 269,  274, 2048+1484,
 275,  280, 2048+1485,
 281,  286, 2048+1486,
 287,  292, 2048+1487,
 293,  298, 2048+1488,
 299,  304, 2048+1489,
 305,  310, 2048+1490,
 311,  316, 2048+1491,
 317,  322, 2048+1492,
 323,  328, 2048+1493,
 329,  334, 2048+1494,
 335,  340, 2048+1495,
 341,  346, 2048+1496,
 347,  352, 2048+1497,
 353,  358, 2048+1498,
 359,  364, 2048+1499,
 365,  370, 2048+1500,
 371,  376, 2048+1501,
 377,  382, 2048+1502,
 383,  388, 2048+1503,
 389,  394, 2048+1504,
 395,  400, 2048+1505,
 401,  406, 2048+1506,
 407,  412, 2048+1507,
 413,  418, 2048+1508,
 419,  424, 2048+1509,
 425,  430, 2048+1510,
 431,  436, 2048+1511,
 437,  442, 2048+1512,
 443,  448, 2048+1513,
 449,  454, 2048+1514,
 455,  460, 2048+1515,
 461,  466, 2048+1516,
 467,  472, 2048+1517,
 473,  478, 2048+1518,
 479,  484, 2048+1519,
 485,  490, 2048+1520,
 491,  496, 2048+1521,
 497,  502, 2048+1522,
 503,  508, 2048+1523,
 509,  514, 2048+1524,
 515,  520, 2048+1525,
 521,  526, 2048+1526,
 527,  532, 2048+1527,
 533,  538, 2048+1528,
 539,  544, 2048+1529,
 545,  550, 2048+1530,
 551,  556, 2048+1531,
 557,  562, 2048+1532,
 563,  568, 2048+1533,
 569,  574, 2048+1534,
 575,  580, 2048+1535,
 581,  586, 2048+1536,
 587,  592, 2048+1537,
 593,  598, 2048+1538,
 599,  604, 2048+1539,
 605,  610, 2048+1540,
 611,  616, 2048+1541,
 617,  622, 2048+1542,
 623,  628, 2048+1543,
 629,  634, 2048+1544,
 635,  640, 2048+1545,
 641,  646, 2048+1546,
 647,  652, 2048+1547,
 653,  658, 2048+1548,
 659,  664, 2048+1549,
 665,  670, 2048+1550,
 671,  676, 2048+1551,
 677,  682, 2048+1552,
 683,  688, 2048+1553,
 689,  694, 2048+1554,
 695,  700, 2048+1555,
 701,  706, 2048+1556,
 707,  712, 2048+1557,
 713,  718, 2048+1558,
 719,  724, 2048+1559,
 725,  730, 2048+1560,
 731,  736, 2048+1561,
 737,  742, 2048+1562,
 743,  748, 2048+1563,
 749,  754, 2048+1564,
 755,  760, 2048+1565,
 761,  766, 2048+1566,
 767,  772, 2048+1567,
 773,  778, 2048+1568,
 779,  784, 2048+1569,
 785,  790, 2048+1570,
 791,  796, 2048+1571,
 797,  802, 2048+1572,
 803,  808, 2048+1573,
 809,  814, 2048+1574,
 815,  820, 2048+1575,
 821,  826, 2048+1576,
 827,  832, 2048+1577,
 833,  838, 2048+1578,
 839,  844, 2048+1579,
 845,  850, 2048+1580,
 851,  856, 2048+1581,
 857,  862, 2048+1582,
 863,  868, 2048+1583,
 869,  874, 2048+1584,
 875,  880, 2048+1585,
 881,  886, 2048+1586,
 887,  892, 2048+1587,
 893,  898, 2048+1588,
 899,  904, 2048+1589,
 905,  910, 2048+1590,
 911,  916, 2048+1591,
 917,  922, 2048+1592,
 923,  928, 2048+1593,
 929,  934, 2048+1594,
 935,  940, 2048+1595,
 941,  946, 2048+1596,
 947,  952, 2048+1597,
 953,  958, 2048+1598,
 959,  964, 2048+1599,
 965,  970, 2048+1600,
 971,  976, 2048+1601,
 977,  982, 2048+1602,
 983,  988, 2048+1603,
 989,  994, 2048+1604,
 995, 1000, 2048+1605,
1001, 1006, 2048+1606,
1007, 1012, 2048+1607,
1013, 1018, 2048+1608,
1019, 1024, 2048+1609,
1025, 1030, 2048+1610,
1031, 1036, 2048+1611,
1037, 1042, 2048+1612,
1043, 1048, 2048+1613,
1049, 1054, 2048+1614,
1055, 1060, 2048+1615,
1061, 1066, 2048+1616,
1067, 1072, 2048+1617,
1073, 1078, 2048+1618,
1079, 1084, 2048+1619,
1085, 1090, 2048+1620,
1091, 1096, 2048+1621,
1097, 1102, 2048+1622,
1103, 1108, 2048+1623,
1109, 1114, 2048+1624,
1115, 1120, 2048+1625,
1121, 1126, 2048+1626,
1127, 1132, 2048+1627,
1133, 1138, 2048+1628,
1139, 1144, 2048+1629,
1145, 1150, 2048+1630,
1151, 1156, 2048+1631,
1157, 1162, 2048+1632,
1163, 1168, 2048+1633,
1169, 1174, 2048+1634,
1175, 1180, 2048+1635,
1181, 1186, 2048+1636,
1187, 1192, 2048+1637,
1193, 1198, 2048+1638,
1199, 1204, 2048+1639,
1205, 1210, 2048+1640,
1211, 1216, 2048+1641,
1217, 1222, 2048+1642,
1223, 1228, 2048+1643,
1229, 1234, 2048+1644,
1235, 1240, 2048+1645,
1241, 1246, 2048+1646,
1247, 1252, 2048+1647,
1253, 1258, 2048+1648,
1259, 1264, 2048+1649,
1265, 1270, 2048+1650,
1271, 1276, 2048+1651,
1277, 1282, 2048+1652,
1283, 1288, 2048+1653,
1289, 1294, 2048+1654,
   5, 1295, 2048+1655,
 834,  840, 1074, 2048+1302,
 378,  438,  756, 2048+1303,
 510,  655, 1284, 2048+1304,
 318,  696, 1044, 2048+1305,
 426,  612,  702, 2048+1306,
 918, 1050, 1224, 2048+1307,
 206,  258, 1164, 2048+1308,
 294,  686,  984, 2048+1309,
 168,  181,  954, 2048+1310,
 300,  714, 1092, 2048+1311,
 835,  924, 1285, 2048+1312,
 324,  409,  546, 2048+1313,
 996, 1002, 1237, 2048+1320,
 541,  600,  919, 2048+1321,
 150,  672,  817, 2048+1322,
 481,  859, 1207, 2048+1323,
 588,  774,  865, 2048+1324,
  90, 1080, 1212, 2048+1325,
  30,  368,  420, 2048+1326,
 456,  849, 1146, 2048+1327,
 331,  343, 1116, 2048+1328,
 462,  876, 1255, 2048+1329,
 151,  997, 1087, 2048+1330,
 486,  571,  708, 2048+1331,
 104, 1158, 1165, 2048+1338,
 704,  762, 1081, 2048+1339,
 312,  836,  979, 2048+1340,
  73,  645, 1021, 2048+1341,
 750,  937, 1027, 2048+1342,
  79,  254, 1242, 2048+1343,
 193,  530,  582, 2048+1344,
  12,  618, 1011, 2048+1345,
 493,  505, 1278, 2048+1346,
 121,  625, 1039, 2048+1347,
 313, 1159, 1250, 2048+1348,
 650,  733,  870, 2048+1349,
  25,   31,  266, 2048+1356,
 867,  925, 1243, 2048+1357,
 475,  998, 1141, 2048+1358,
 237,  807, 1183, 2048+1359,
 912, 1100, 1189, 2048+1360,
 109,  241,  416, 2048+1361,
 355,  692,  744, 2048+1362,
 174,  781, 1173, 2048+1363,
 147,  657,  667, 2048+1364,
 284,  787, 1202, 2048+1365,
  26,  116,  476, 2048+1366,
 812,  895, 1033, 2048+1367,
 187,  194,  429, 2048+1374,
 110, 1029, 1088, 2048+1375,
   7,  637, 1160, 2048+1376,
  49,  399,  969, 2048+1377,
  55, 1075, 1262, 2048+1378,
 271,  404,  578, 2048+1379,
 517,  855,  907, 2048+1380,
  39,  336,  943, 2048+1381,
 309,  819,  830, 2048+1382,
  69,  447,  950, 2048+1383,
 188,  278,  638, 2048+1384,
 974, 1057, 1196, 2048+1385,
 349,  356,  591, 2048+1392,
 272, 1191, 1251, 2048+1393,
  27,  170,  799, 2048+1394,
 212,  561, 1131, 2048+1395,
 128,  217, 1238, 2048+1396,
 434,  567,  741, 2048+1397,
 680, 1017, 1070, 2048+1398,
 201,  499, 1105, 2048+1399,
 471,  981,  992, 2048+1400,
 231,  609, 1112, 2048+1401,
 350,  441,  800, 2048+1402,
  63, 1137, 1221, 2048+1403,
 512,  518,  753, 2048+1410,
  57,  117,  435, 2048+1411,
 189,  333,  961, 2048+1412,
 374,  723, 1293, 2048+1413,
 105,  291,  380, 2048+1414,
 596,  729,  903, 2048+1415,
 843, 1179, 1232, 2048+1416,
 363,  663, 1267, 2048+1417,
 633, 1143, 1154, 2048+1418,
 393,  771, 1275, 2048+1419,
 513,  603,  962, 2048+1420,
   3,   87,  225, 2048+1421,
 674,  681,  915, 2048+1428,
 219,  279,  597, 2048+1429,
 351,  495, 1124, 2048+1430,
 159,  537,  885, 2048+1431,
 267,  453,  543, 2048+1432,
 759,  891, 1065, 2048+1433,
  45,   99, 1005, 2048+1434,
 135,  525,  825, 2048+1435,
   9,   21,  795, 2048+1436,
 141,  555,  933, 2048+1437,
 675,  765, 1125, 2048+1438,
 165,  249,  387, 2048+1439,
  60,  144,  204,  234,  235,  288,  474,  540,  660,  906, 1068, 1218, 2048+1296,
  18,   78,  145,  252,  330,  480,  642, 1038, 1098, 1194, 1248, 1254, 2048+1297,
  96,  132,  180,  444,  534,  624,  684,  738,  780,  828, 1206, 1219, 2048+1298,
  24,  102,  108,  205,  210,  564,  648,  654,  685, 1122, 1236, 1272, 2048+1299,
  66,  133,  146,  192,  282,  643,  649,  678,  846,  858,  936, 1086, 2048+1300,
 253,  402,  408,  432,  498,  661,  852,  864,  948, 1032, 1134, 1200, 2048+1301,
  84,  222,  306,  366,  396,  397,  450,  636,  703,  822, 1069, 1230, 2048+1314,
  61,  114,  120,  182,  240,  307,  414,  492,  644,  804, 1201, 1260, 2048+1315,
  72,   85,  259,  295,  342,  606,  697,  786,  847,  900,  942,  990, 2048+1316,
 103,  138,  186,  264,  270,  367,  372,  726,  810,  816,  848, 1286, 2048+1317,
 228,  296,  308,  354,  445,  805,  811,  841, 1008, 1020, 1099, 1249, 2048+1318,
   0,   67,  415,  565,  570,  594,  662,  823, 1014, 1026, 1110, 1195, 2048+1319,
  97,  246,  384,  468,  528,  558,  559,  613,  798,  866,  985, 1231, 2048+1332,
  68,  126,  223,  276,  283,  344,  403,  469,  576,  656,  806,  966, 2048+1333,
 236,  247,  421,  457,  504,  768,  860,  949, 1009, 1062, 1104, 1152, 2048+1334,
 152,  265,  301,  348,  427,  433,  529,  535,  888,  972,  978, 1010, 2048+1335,
 115,  390,  458,  470,  516,  607,  967,  973, 1003, 1170, 1182, 1261, 2048+1336,
  62,  162,  229,  577,  727,  732,  757,  824,  986, 1176, 1188, 1273, 2048+1337,
  98,  260,  410,  547,  630,  690,  720,  721,  775,  960, 1028, 1147, 2048+1350,
 230,  289,  385,  439,  446,  506,  566,  631,  739,  818,  968, 1128, 2048+1351,
  19,  398,  411,  583,  619,  666,  930, 1022, 1111, 1171, 1225, 1266, 2048+1352,
 314,  428,  463,  511,  589,  595,  691,  698, 1051, 1135, 1140, 1172, 2048+1353,
  36,   48,  127,  277,  552,  620,  632,  679,  769, 1129, 1136, 1166, 2048+1354,
  42,   54,  139,  224,  325,  391,  740,  889,  894,  920,  987, 1148, 2048+1355,
  13,  261,  422,  572,  709,  792,  853,  882,  883,  938, 1123, 1190, 2048+1368,
 392,  451,  548,  601,  608,  668,  728,  793,  901,  980, 1130, 1290, 2048+1369,
  37,   91,  134,  183,  560,  573,  745,  782,  829, 1093, 1184, 1274, 2048+1370,
   1,    6,   38,  477,  590,  626,  673,  751,  758,  854,  861, 1213, 2048+1371,
   2,   32,  198,  211,  290,  440,  715,  783,  794,  842,  931, 1291, 2048+1372,
  14,  207,  216,  302,  386,  487,  553,  902, 1052, 1056, 1082, 1149, 2048+1373,
  56,  175,  423,  584,  734,  871,  955, 1015, 1045, 1046, 1101, 1287, 2048+1386,
 156,  554,  614,  710,  763,  770,  831,  890,  956, 1063, 1142, 1292, 2048+1387,
  50,  140,  199,  255,  297,  345,  722,  735,  908,  944,  991, 1256, 2048+1388,
  80,  163,  169,  200,  639,  752,  788,  837,  913,  921, 1016, 1023, 2048+1389,
 157,  164,  195,  360,  373,  452,  602,  877,  945,  957, 1004, 1094, 2048+1390,
  15,  176,  369,  379,  464,  549,  651,  716, 1064, 1214, 1220, 1244, 2048+1391,
 153,  218,  337,  585,  746,  896, 1034, 1117, 1177, 1208, 1209, 1263, 2048+1404,
   8,  158,  319,  717,  776,  872,  926,  932,  993, 1053, 1118, 1226, 2048+1405,
 122,  213,  303,  361,  417,  459,  507,  884,  897, 1071, 1106, 1153, 2048+1406,
 242,  326,  332,  362,  801,  914,  951,  999, 1076, 1083, 1178, 1185, 2048+1407,
 320,  327,  357,  522,  536,  615,  764, 1040, 1107, 1119, 1167, 1257, 2048+1408,
  81,   86,  111,  177,  338,  531,  542,  627,  711,  813,  878, 1227, 2048+1409,
  43,   74,   75,  129,  315,  381,  500,  747,  909, 1058, 1197, 1279, 2048+1422,
  92,  171,  321,  482,  879,  939, 1035, 1089, 1095, 1155, 1215, 1280, 2048+1423,
  20,  285,  375,  465,  523,  579,  621,  669, 1047, 1059, 1233, 1268, 2048+1424,
  44,   51,  405,  488,  494,  524,  963, 1077, 1113, 1161, 1239, 1245, 2048+1425,
  33,  123,  483,  489,  519,  687,  699,  777,  927, 1203, 1269, 1281, 2048+1426,
  93,  243,  248,  273,  339,  501,  693,  705,  789,  873,  975, 1041, 2048+1427,

   3,    9, 2048+1240,
  10,   16, 2048+1241,
  17,   22, 2048+1242,
  23,   26, 2048+1243,
  27,   31, 2048+1244,
  32,   35, 2048+1245,
  36,   40, 2048+1246,
  41,   46, 2048+1247,
  47,   51, 2048+1248,
  52,   56, 2048+1249,
  57,   62, 2048+1250,
  63,   68, 2048+1251,
  69,   74, 2048+1252,
  75,   80, 2048+1253,
  81,   85, 2048+1254,
  86,   89, 2048+1255,
  90,   95, 2048+1256,
  96,  100, 2048+1257,
 101,  104, 2048+1258,
 105,  110, 2048+1259,
 111,  115, 2048+1260,
 116,  121, 2048+1261,
 122,  126, 2048+1262,
 127,  133, 2048+1263,
 134,  138, 2048+1264,
 139,  144, 2048+1265,
 145,  151, 2048+1266,
 152,  157, 2048+1267,
 158,  161, 2048+1268,
 162,  166, 2048+1269,
 167,  170, 2048+1270,
 171,  175, 2048+1271,
 176,  181, 2048+1272,
 182,  186, 2048+1273,
 187,  191, 2048+1274,
 192,  197, 2048+1275,
 198,  203, 2048+1276,
 204,  209, 2048+1277,
 210,  215, 2048+1278,
 216,  220, 2048+1279,
 221,  224, 2048+1280,
 225,  230, 2048+1281,
 231,  235, 2048+1282,
 236,  239, 2048+1283,
 240,  245, 2048+1284,
 246,  250, 2048+1285,
 251,  256, 2048+1286,
 257,  261, 2048+1287,
 262,  268, 2048+1288,
 269,  273, 2048+1289,
 274,  279, 2048+1290,
 280,  286, 2048+1291,
 287,  292, 2048+1292,
 293,  296, 2048+1293,
 297,  301, 2048+1294,
 302,  305, 2048+1295,
 306,  310, 2048+1296,
 311,  316, 2048+1297,
 317,  321, 2048+1298,
 322,  326, 2048+1299,
 327,  332, 2048+1300,
 333,  338, 2048+1301,
 339,  344, 2048+1302,
 345,  350, 2048+1303,
 351,  355, 2048+1304,
 356,  359, 2048+1305,
 360,  365, 2048+1306,
 366,  370, 2048+1307,
 371,  374, 2048+1308,
 375,  380, 2048+1309,
 381,  385, 2048+1310,
 386,  391, 2048+1311,
 392,  396, 2048+1312,
 397,  403, 2048+1313,
 404,  408, 2048+1314,
 409,  414, 2048+1315,
 415,  421, 2048+1316,
 422,  427, 2048+1317,
 428,  431, 2048+1318,
 432,  436, 2048+1319,
 437,  440, 2048+1320,
 441,  445, 2048+1321,
 446,  451, 2048+1322,
 452,  456, 2048+1323,
 457,  461, 2048+1324,
 462,  467, 2048+1325,
 468,  473, 2048+1326,
 474,  479, 2048+1327,
 480,  485, 2048+1328,
 486,  490, 2048+1329,
 491,  494, 2048+1330,
 495,  500, 2048+1331,
 501,  505, 2048+1332,
 506,  509, 2048+1333,
 510,  515, 2048+1334,
 516,  520, 2048+1335,
 521,  526, 2048+1336,
 527,  531, 2048+1337,
 532,  538, 2048+1338,
 539,  543, 2048+1339,
 544,  549, 2048+1340,
 550,  556, 2048+1341,
 557,  562, 2048+1342,
 563,  566, 2048+1343,
 567,  571, 2048+1344,
 572,  575, 2048+1345,
 576,  580, 2048+1346,
 581,  586, 2048+1347,
 587,  591, 2048+1348,
 592,  596, 2048+1349,
 597,  602, 2048+1350,
 603,  608, 2048+1351,
 609,  614, 2048+1352,
 615,  620, 2048+1353,
 621,  625, 2048+1354,
 626,  629, 2048+1355,
 630,  635, 2048+1356,
 636,  640, 2048+1357,
 641,  644, 2048+1358,
 645,  650, 2048+1359,
 651,  655, 2048+1360,
 656,  661, 2048+1361,
 662,  666, 2048+1362,
 667,  673, 2048+1363,
 674,  678, 2048+1364,
 679,  684, 2048+1365,
 685,  691, 2048+1366,
 692,  697, 2048+1367,
 698,  701, 2048+1368,
 702,  706, 2048+1369,
 707,  710, 2048+1370,
 711,  715, 2048+1371,
 716,  721, 2048+1372,
 722,  726, 2048+1373,
 727,  731, 2048+1374,
 732,  737, 2048+1375,
 738,  743, 2048+1376,
 744,  749, 2048+1377,
 750,  755, 2048+1378,
 756,  760, 2048+1379,
 761,  764, 2048+1380,
 765,  770, 2048+1381,
 771,  775, 2048+1382,
 776,  779, 2048+1383,
 780,  785, 2048+1384,
 786,  790, 2048+1385,
 791,  796, 2048+1386,
 797,  801, 2048+1387,
 802,  808, 2048+1388,
 809,  813, 2048+1389,
 814,  819, 2048+1390,
 820,  826, 2048+1391,
 827,  832, 2048+1392,
 833,  836, 2048+1393,
 837,  841, 2048+1394,
 842,  845, 2048+1395,
 846,  850, 2048+1396,
 851,  856, 2048+1397,
 857,  861, 2048+1398,
 862,  866, 2048+1399,
 867,  872, 2048+1400,
 873,  878, 2048+1401,
 879,  884, 2048+1402,
 885,  890, 2048+1403,
 891,  895, 2048+1404,
 896,  899, 2048+1405,
 900,  905, 2048+1406,
 906,  910, 2048+1407,
 911,  914, 2048+1408,
 915,  920, 2048+1409,
 921,  925, 2048+1410,
 926,  931, 2048+1411,
 932,  936, 2048+1412,
 937,  943, 2048+1413,
 944,  948, 2048+1414,
 949,  954, 2048+1415,
 955,  961, 2048+1416,
 962,  967, 2048+1417,
 968,  971, 2048+1418,
 972,  976, 2048+1419,
 977,  980, 2048+1420,
 981,  985, 2048+1421,
 986,  991, 2048+1422,
 992,  996, 2048+1423,
 997, 1001, 2048+1424,
1002, 1007, 2048+1425,
1008, 1013, 2048+1426,
1014, 1019, 2048+1427,
1020, 1025, 2048+1428,
1026, 1030, 2048+1429,
1031, 1034, 2048+1430,
1035, 1040, 2048+1431,
1041, 1045, 2048+1432,
1046, 1049, 2048+1433,
1050, 1055, 2048+1434,
1056, 1060, 2048+1435,
1061, 1066, 2048+1436,
1067, 1071, 2048+1437,
1072, 1078, 2048+1438,
   4, 1079, 2048+1439,
   0,  247,  723, 2048+1085,
   5,  298,  357, 2048+1086,
  13,   64,  507, 2048+1087,
  19,  211,  853, 2048+1088,
  24,  119,  270, 2048+1089,
  28,  487,  669, 2048+1090,
  33,  264,  362, 2048+1091,
  37,  107,  226, 2048+1092,
  34,   42,  433, 2048+1093,
  48,  177,  416, 2048+1094,
  53,  367,  453, 2048+1095,
  58,  728, 1057, 2048+1096,
  65,  153,  886, 2048+1097,
  70,  307, 1015, 2048+1098,
  59,   76,  271, 2048+1099,
 135,  382,  858, 2048+1105,
 140,  434,  493, 2048+1106,
 148,  199,  642, 2048+1107,
 155,  346,  988, 2048+1108,
 159,  254,  405, 2048+1109,
 163,  622,  804, 2048+1110,
 168,  399,  497, 2048+1111,
 172,  243,  363, 2048+1112,
 169,  178,  568, 2048+1113,
 183,  312,  551, 2048+1114,
 188,  503,  588, 2048+1115,
 113,  193,  863, 2048+1116,
 200,  288, 1021, 2048+1117,
  71,  206,  442, 2048+1118,
 194,  212,  406, 2048+1119,
 272,  517,  993, 2048+1125,
 275,  569,  628, 2048+1126,
 283,  335,  777, 2048+1127,
  44,  290,  482, 2048+1128,
 294,  389,  540, 2048+1129,
 299,  758,  939, 2048+1130,
 303,  534,  632, 2048+1131,
 308,  378,  498, 2048+1132,
 304,  313,  703, 2048+1133,
 318,  447,  686, 2048+1134,
 323,  638,  724, 2048+1135,
 249,  329,  999, 2048+1136,
  77,  336,  423, 2048+1137,
 207,  342,  578, 2048+1138,
 330,  347,  541, 2048+1139,
  49,  407,  652, 2048+1145,
 411,  704,  763, 2048+1146,
 419,  470,  912, 2048+1147,
 180,  425,  617, 2048+1148,
 429,  525,  675, 2048+1149,
 435,  893, 1074, 2048+1150,
 438,  671,  768, 2048+1151,
 443,  513,  633, 2048+1152,
 439,  448,  838, 2048+1153,
 454,  582,  821, 2048+1154,
 458,  774,  859, 2048+1155,
  55,  384,  464, 2048+1156,
 213,  471,  558, 2048+1157,
 343,  477,  713, 2048+1158,
 465,  483,  676, 2048+1159,
 184,  542,  787, 2048+1165,
 547,  839,  898, 2048+1166,
 554,  606, 1047, 2048+1167,
 315,  560,  752, 2048+1168,
 564,  660,  810, 2048+1169,
 130,  570, 1029, 2048+1170,
 573,  806,  903, 2048+1171,
 579,  649,  769, 2048+1172,
 574,  583,  973, 2048+1173,
 589,  717,  957, 2048+1174,
 593,  909,  994, 2048+1175,
 190,  519,  599, 2048+1176,
 348,  607,  694, 2048+1177,
 478,  612,  848, 2048+1178,
 600,  618,  811, 2048+1179,
 319,  677,  922, 2048+1185,
 683,  974, 1033, 2048+1186,
 102,  689,  741, 2048+1187,
 450,  696,  888, 2048+1188,
 699,  795,  945, 2048+1189,
  84,  267,  705, 2048+1190,
 708,  941, 1038, 2048+1191,
 714,  784,  904, 2048+1192,
  29,  709,  718, 2048+1193,
  15,  725,  854, 2048+1194,
  50,  729, 1044, 2048+1195,
 325,  654,  734, 2048+1196,
 484,  742,  829, 2048+1197,
 613,  747,  983, 2048+1198,
 735,  753,  946, 2048+1199,
 455,  812, 1058, 2048+1205,
  30,   88,  818, 2048+1206,
 237,  824,  876, 2048+1207,
 585,  831, 1023, 2048+1208,
   1,  835,  930, 2048+1209,
 219,  402,  840, 2048+1210,
  93,  843, 1076, 2048+1211,
 849,  919, 1039, 2048+1212,
 164,  844,  855, 2048+1213,
 150,  860,  989, 2048+1214,
  99,  185,  864, 2048+1215,
 460,  789,  869, 2048+1216,
 619,  877,  964, 2048+1217,
  39,  748,  882, 2048+1218,
   2,  870,  889, 2048+1219,
 114,  590,  947, 2048+1225,
 165,  223,  953, 2048+1226,
 373,  960, 1011, 2048+1227,
  79,  720,  966, 2048+1228,
 136,  970, 1065, 2048+1229,
 354,  537,  975, 2048+1230,
 132,  229,  978, 2048+1231,
  94,  984, 1054, 2048+1232,
 300,  979,  990, 2048+1233,
  45,  285,  995, 2048+1234,
 234,  320, 1000, 2048+1235,
 595,  924, 1005, 2048+1236,
  21,  754, 1012, 2048+1237,
 174,  883, 1018, 2048+1238,
 137, 1006, 1024, 2048+1239,
 106,  241,  328,  334,  604,  834,  852, 1003, 2048+1080,
 112,  117,  410,  481,  693,  772,  798,  799, 2048+1081,
 118,  205,  372,  502,  545,  577,  680, 1027, 2048+1082,
  11,  123,  263,  361,  492,  646,  668,  956, 2048+1083,
  12,   18,  128,  340,  522,  757,  766,  998, 2048+1084,
  60,  242,  376,  463,  469,  739,  969,  987, 2048+1100,
 248,  252,  546,  616,  828,  907,  933,  934, 2048+1101,
  82,  253,  341,  508,  637,  681,  712,  815, 2048+1102,
  14,  146,  258,  398,  496,  627,  781,  803, 2048+1103,
  54,  147,  154,  265,  475,  657,  892,  901, 2048+1104,
  25,   43,  195,  377,  511,  598,  605,  874, 2048+1120,
 383,  387,  682,  751,  963, 1042, 1068, 1069, 2048+1121,
 217,  388,  476,  643,  773,  816,  847,  950, 2048+1122,
 149,  281,  393,  533,  631,  762,  916,  938, 2048+1123,
 189,  282,  289,  400,  610,  792, 1028, 1036, 2048+1124,
 160,  179,  331,  512,  647,  733,  740, 1009, 2048+1140,
  20,   97,  124,  125,  518,  523,  817,  887, 2048+1141,
   6,  352,  524,  611,  778,  908,  951,  982, 2048+1142,
 284,  417,  528,  670,  767,  897, 1051, 1073, 2048+1143,
  83,   91,  324,  418,  424,  535,  745,  927, 2048+1144,
  66,  295,  314,  466,  648,  782,  868,  875, 2048+1160,
 156,  232,  259,  260,  653,  658,  952, 1022, 2048+1161,
   7,   38,  141,  488,  659,  746,  913, 1043, 2048+1162,
 108,  129,  420,  552,  663,  805,  902, 1032, 2048+1163,
 218,  227,  459,  553,  559,  672,  880, 1062, 2048+1164,
 201,  430,  449,  601,  783,  917, 1004, 1010, 2048+1180,
   8,   78,  291,  368,  394,  395,  788,  793, 2048+1181,
  98,  142,  173,  276,  623,  794,  881, 1048, 2048+1182,
  87,  244,  266,  555,  687,  800,  940, 1037, 2048+1183,
 120,  353,  364,  594,  688,  695,  807, 1016, 2048+1184,
  61,   67,  337,  565,  584,  736,  918, 1052, 2048+1200,
 143,  214,  426,  504,  529,  530,  923,  928, 2048+1201,
 103,  233,  277,  309,  412,  759,  929, 1017, 2048+1202,
  92,  222,  379,  401,  690,  822,  935, 1075, 2048+1203,
  72,  255,  489,  499,  730,  823,  830,  942, 2048+1204,
 109,  196,  202,  472,  700,  719,  871, 1053, 2048+1220,
 278,  349,  561,  639,  664,  665, 1059, 1063, 2048+1221,
  73,  238,  369,  413,  444,  548,  894, 1064, 2048+1222,
 131,  228,  358,  514,  536,  825,  958, 1070, 2048+1223,
 208,  390,  624,  634,  865,  959,  965, 1077, 2048+1224,

   9,   20, 2048+1800,
  21,   31, 2048+1801,
  32,   42, 2048+1802,
  43,   53, 2048+1803,
  54,   64, 2048+1804,
  65,   75, 2048+1805,
  76,   86, 2048+1806,
  87,   97, 2048+1807,
  98,  108, 2048+1808,
 109,  119, 2048+1809,
 120,  130, 2048+1810,
 131,  141, 2048+1811,
 142,  152, 2048+1812,
 153,  163, 2048+1813,
 164,  174, 2048+1814,
 175,  185, 2048+1815,
 186,  196, 2048+1816,
 197,  207, 2048+1817,
 208,  218, 2048+1818,
 219,  229, 2048+1819,
 230,  240, 2048+1820,
 241,  251, 2048+1821,
 252,  262, 2048+1822,
 263,  273, 2048+1823,
 274,  284, 2048+1824,
 285,  295, 2048+1825,
 296,  306, 2048+1826,
 307,  317, 2048+1827,
 318,  328, 2048+1828,
 329,  339, 2048+1829,
 340,  350, 2048+1830,
 351,  361, 2048+1831,
 362,  372, 2048+1832,
 373,  383, 2048+1833,
 384,  394, 2048+1834,
 395,  405, 2048+1835,
 406,  416, 2048+1836,
 417,  427, 2048+1837,
 428,  438, 2048+1838,
 439,  449, 2048+1839,
 450,  460, 2048+1840,
 461,  471, 2048+1841,
 472,  482, 2048+1842,
 483,  493, 2048+1843,
 494,  504, 2048+1844,
 505,  515, 2048+1845,
 516,  526, 2048+1846,
 527,  537, 2048+1847,
 538,  548, 2048+1848,
 549,  559, 2048+1849,
 560,  570, 2048+1850,
 571,  581, 2048+1851,
 582,  592, 2048+1852,
 593,  603, 2048+1853,
 604,  614, 2048+1854,
 615,  625, 2048+1855,
 626,  636, 2048+1856,
 637,  647, 2048+1857,
 648,  658, 2048+1858,
 659,  669, 2048+1859,
 670,  680, 2048+1860,
 681,  691, 2048+1861,
 692,  702, 2048+1862,
 703,  713, 2048+1863,
 714,  724, 2048+1864,
 725,  735, 2048+1865,
 736,  746, 2048+1866,
 747,  757, 2048+1867,
 758,  768, 2048+1868,
 769,  779, 2048+1869,
 780,  790, 2048+1870,
 791,  801, 2048+1871,
 802,  812, 2048+1872,
 813,  823, 2048+1873,
 824,  834, 2048+1874,
 835,  845, 2048+1875,
 846,  856, 2048+1876,
 857,  867, 2048+1877,
 868,  878, 2048+1878,
 879,  889, 2048+1879,
 890,  900, 2048+1880,
 901,  911, 2048+1881,
 912,  922, 2048+1882,
 923,  933, 2048+1883,
 934,  944, 2048+1884,
 945,  955, 2048+1885,
 956,  966, 2048+1886,
 967,  977, 2048+1887,
 978,  988, 2048+1888,
 989,  999, 2048+1889,
1000, 1010, 2048+1890,
1011, 1021, 2048+1891,
1022, 1032, 2048+1892,
1033, 1043, 2048+1893,
1044, 1054, 2048+1894,
1055, 1065, 2048+1895,
1066, 1076, 2048+1896,
1077, 1087, 2048+1897,
1088, 1098, 2048+1898,
1099, 1109, 2048+1899,
1110, 1120, 2048+1900,
1121, 1131, 2048+1901,
1132, 1142, 2048+1902,
1143, 1153, 2048+1903,
1154, 1164, 2048+1904,
1165, 1175, 2048+1905,
1176, 1186, 2048+1906,
1187, 1197, 2048+1907,
1198, 1208, 2048+1908,
1209, 1219, 2048+1909,
1220, 1230, 2048+1910,
1231, 1241, 2048+1911,
1242, 1252, 2048+1912,
1253, 1263, 2048+1913,
1264, 1274, 2048+1914,
1275, 1285, 2048+1915,
1286, 1296, 2048+1916,
1297, 1307, 2048+1917,
1308, 1318, 2048+1918,
1319, 1329, 2048+1919,
1330, 1340, 2048+1920,
1341, 1351, 2048+1921,
1352, 1362, 2048+1922,
1363, 1373, 2048+1923,
1374, 1384, 2048+1924,
1385, 1395, 2048+1925,
1396, 1406, 2048+1926,
1407, 1417, 2048+1927,
1418, 1428, 2048+1928,
1429, 1439, 2048+1929,
1440, 1450, 2048+1930,
1451, 1461, 2048+1931,
1462, 1472, 2048+1932,
1473, 1483, 2048+1933,
1484, 1494, 2048+1934,
1495, 1505, 2048+1935,
1506, 1516, 2048+1936,
1517, 1527, 2048+1937,
1528, 1538, 2048+1938,
1539, 1549, 2048+1939,
1550, 1560, 2048+1940,
1561, 1571, 2048+1941,
1572, 1582, 2048+1942,
  10, 1583, 2048+1943,
   0,   11,  671, 2048+1593,
  12,  231,  924, 2048+1594,
  22,  594, 1177, 2048+1595,
  35,  540,  913, 2048+1596,
  44,  154,  892, 2048+1597,
  56,   57, 1366, 2048+1598,
  66,  463,  704, 2048+1599,
  78, 1012, 1276, 2048+1600,
  88,  836, 1156, 2048+1601,
  99, 1343, 1387, 2048+1602,
 111,  188,  869, 2048+1603,
 122,  123,  541, 2048+1604,
 132,  254, 1476, 2048+1605,
 143,  429, 1299, 2048+1606,
 155,  265, 1090, 2048+1607,
 165,  572,  837, 2048+1608,
 177,  759, 1013, 2048+1609,
  13,  133,  189, 2048+1610,
 198,  209,  870, 2048+1620,
 210,  430, 1122, 2048+1621,
 221,  794, 1375, 2048+1622,
 234,  739, 1111, 2048+1623,
 243,  352, 1092, 2048+1624,
 256,  257, 1565, 2048+1625,
 266,  662,  903, 2048+1626,
 277, 1211, 1477, 2048+1627,
 288, 1036, 1355, 2048+1628,
   2,  297, 1543, 2048+1629,
 309,  386, 1069, 2048+1630,
 322,  323,  740, 2048+1631,
  91,  330,  452, 2048+1632,
 342,  628, 1498, 2048+1633,
 353,  465, 1290, 2048+1634,
 363,  771, 1037, 2048+1635,
 375,  959, 1212, 2048+1636,
 211,  331,  387, 2048+1637,
 396,  409, 1070, 2048+1647,
 410,  629, 1321, 2048+1648,
 421,  993, 1575, 2048+1649,
 433,  937, 1309, 2048+1650,
 441,  550, 1292, 2048+1651,
 181,  454,  455, 2048+1652,
 466,  862, 1102, 2048+1653,
  92,  476, 1411, 2048+1654,
 487, 1235, 1554, 2048+1655,
 159,  200,  495, 2048+1656,
 508,  585, 1267, 2048+1657,
 521,  522,  938, 2048+1658,
 291,  532,  652, 2048+1659,
 114,  543,  826, 2048+1660,
 551,  664, 1489, 2048+1661,
 562,  969, 1236, 2048+1662,
 574, 1159, 1412, 2048+1663,
 411,  533,  586, 2048+1664,
 595,  608, 1268, 2048+1674,
 609,  827, 1519, 2048+1675,
 192,  619, 1193, 2048+1676,
 632, 1135, 1509, 2048+1677,
 640,  750, 1491, 2048+1678,
 379,  654,  655, 2048+1679,
 665, 1060, 1302, 2048+1680,
  26,  292,  675, 2048+1681,
 169,  686, 1434, 2048+1682,
 357,  398,  694, 2048+1683,
 707,  784, 1466, 2048+1684,
 719,  720, 1136, 2048+1685,
 490,  731,  850, 2048+1686,
 312,  742, 1024, 2048+1687,
 104,  751,  864, 2048+1688,
 761, 1168, 1435, 2048+1689,
  27,  773, 1358, 2048+1690,
 610,  732,  785, 2048+1691,
 795,  807, 1467, 2048+1701,
 135,  808, 1025, 2048+1702,
 390,  817, 1393, 2048+1703,
 126,  830, 1335, 2048+1704,
 106,  840,  948, 2048+1705,
 578,  852,  853, 2048+1706,
 865, 1259, 1501, 2048+1707,
 225,  491,  874, 2048+1708,
  49,  367,  884, 2048+1709,
 555,  597,  894, 2048+1710,
  82,  906,  983, 2048+1711,
 918,  919, 1336, 2048+1712,
 689,  930, 1048, 2048+1713,
 511,  940, 1223, 2048+1714,
 302,  949, 1062, 2048+1715,
  50,  961, 1369, 2048+1716,
 226,  971, 1557, 2048+1717,
 809,  931,  984, 2048+1718,
  83,  994, 1005, 2048+1728,
 333, 1006, 1224, 2048+1729,
   8,  589, 1017, 2048+1730,
 326, 1028, 1534, 2048+1731,
 304, 1040, 1147, 2048+1732,
 777, 1050, 1051, 2048+1733,
 117, 1063, 1457, 2048+1734,
 425,  690, 1074, 2048+1735,
 248,  566, 1082, 2048+1736,
 755,  797, 1094, 2048+1737,
 281, 1105, 1182, 2048+1738,
1116, 1117, 1535, 2048+1739,
 887, 1128, 1247, 2048+1740,
 710, 1138, 1423, 2048+1741,
 500, 1148, 1261, 2048+1742,
 249, 1161, 1568, 2048+1743,
 172,  426, 1170, 2048+1744,
1007, 1129, 1183, 2048+1745,
 282, 1194, 1203, 2048+1755,
 535, 1204, 1424, 2048+1756,
 206,  788, 1216, 2048+1757,
 149,  525, 1227, 2048+1758,
 502, 1239, 1347, 2048+1759,
 975, 1249, 1250, 2048+1760,
  72,  315, 1262, 2048+1761,
 623,  888, 1272, 2048+1762,
 446,  765, 1281, 2048+1763,
 953,  996, 1294, 2048+1764,
 480, 1305, 1380, 2048+1765,
 150, 1314, 1315, 2048+1766,
1085, 1327, 1446, 2048+1767,
  40,  909, 1338, 2048+1768,
 699, 1348, 1459, 2048+1769,
 184,  447, 1360, 2048+1770,
 370,  624, 1371, 2048+1771,
1205, 1328, 1381, 2048+1772,
 481, 1394, 1403, 2048+1782,
  41,  734, 1404, 2048+1783,
 404,  987, 1416, 2048+1784,
 348,  723, 1427, 2048+1785,
 701, 1438, 1547, 2048+1786,
1174, 1448, 1449, 2048+1787,
 272,  514, 1460, 2048+1788,
 821, 1086, 1471, 2048+1789,
 645,  965, 1482, 2048+1790,
1152, 1196, 1493, 2048+1791,
 679, 1504, 1580, 2048+1792,
 349, 1514, 1515, 2048+1793,
  63, 1284, 1525, 2048+1794,
 239, 1108, 1537, 2048+1795,
  74,  899, 1548, 2048+1796,
 382,  646, 1559, 2048+1797,
 569,  822, 1570, 2048+1798,
1405, 1526, 1581, 2048+1799,
 242,  319,  561,  649,  858,  902,  990, 1067, 1144, 1232, 1474, 1540, 2048+1584,
  33,  253,  528,  529,  605,  737,  979, 1034, 1210, 1331, 1353, 1419, 2048+1585,
 187,  473,  506,  726,  792, 1166, 1221, 1254, 1342, 1397, 1408, 1409, 2048+1586,
  55,  517,  530,  748, 1100, 1188, 1441, 1463, 1485, 1507, 1551, 1562, 2048+1587,
  34,  110,  176,  275,  650,  693,  803, 1287, 1364, 1365, 1508, 1541, 2048+1588,
 462,  531,  539,  627,  682,  770,  859,  891, 1089, 1398, 1420, 1496, 2048+1589,
  77,  121,  286,  407,  418,  484,  583,  793,  957, 1068, 1155, 1288, 2048+1590,
 264,  287,  320,  749,  958, 1243, 1298, 1320, 1332, 1475, 1529, 1573, 2048+1591,
 220,  341,  408,  419,  638,  660,  781, 1035, 1189, 1386, 1430, 1574, 2048+1592,
  89,  156,  440,  518,  760,  847, 1056, 1101, 1190, 1265, 1344, 1431, 2048+1611,
  36,  232,  451,  727,  728,  804,  935, 1178, 1233, 1410, 1530, 1552, 2048+1612,
  14,   23,   24,  385,  672,  705,  925,  991, 1367, 1421, 1452, 1542, 2048+1613,
  58,   79,  100,  124,  166,  178,  255,  715,  729,  946, 1300, 1388, 2048+1614,
 125,  157,  233,  308,  374,  474,  848,  893, 1001, 1486, 1563, 1564, 2048+1615,
  15,   37,  112,  661,  730,  738,  825,  880,  968, 1057, 1091, 1289, 2048+1616,
 276,  321,  485,  606,  616,  683,  782,  992, 1157, 1266, 1354, 1487, 2048+1617,
  90,  144,  190,  464,  486,  519,  947, 1158, 1442, 1497, 1518, 1531, 2048+1618,
   1,   45,  191,  420,  542,  607,  617,  838,  860,  980, 1234, 1389, 2048+1619,
  46,  289,  354,  639,  716,  960, 1045, 1255, 1301, 1390, 1464, 1544, 2048+1638,
  25,  145,  167,  235,  431,  651,  926,  927, 1002, 1133, 1376, 1432, 2048+1639,
  38,   67,  158,  212,  222,  223,  584,  871,  904, 1123, 1191, 1566, 2048+1640,
   3,  258,  278,  298,  324,  364,  376,  453,  914,  928, 1145, 1499, 2048+1641,
 101,  179,  180,  325,  355,  432,  507,  573,  673, 1046, 1093, 1199, 2048+1642,
 213,  236,  310,  861,  929,  936, 1023, 1078, 1167, 1256, 1291, 1488, 2048+1643,
 102,  475,  520,  684,  805,  814,  881,  981, 1192, 1356, 1465, 1553, 2048+1644,
  59,  113,  134,  146,  290,  343,  388,  663,  685,  717, 1146, 1357, 2048+1645,
   4,  199,  244,  389,  618,  741,  806,  815, 1038, 1058, 1179, 1433, 2048+1646,
   5,   80,  160,  245,  488,  552,  839,  915, 1160, 1244, 1453, 1500, 2048+1665,
  47,  224,  344,  365,  434,  630,  849, 1124, 1125, 1200, 1333, 1576, 2048+1666,
 182,  237,  267,  356,  412,  422,  423,  783, 1071, 1103, 1322, 1391, 2048+1667,
 115,  201,  456,  477,  496,  523,  563,  575,  653, 1112, 1126, 1345, 2048+1668,
 299,  377,  378,  524,  553,  631,  706,  772,  872, 1245, 1293, 1399, 2048+1669,
 103,  413,  435,  509, 1059, 1127, 1134, 1222, 1277, 1368, 1454, 1490, 2048+1670,
  81,  168,  300,  674,  718,  882, 1003, 1014, 1079, 1180, 1392, 1555, 2048+1671,
 259,  311,  332,  345,  489,  544,  587,  863,  883,  916, 1346, 1556, 2048+1672,
  48,  202,  397,  442,  588,  816,  939, 1004, 1015, 1237, 1257, 1377, 2048+1673,
  68,  116,  203,  279,  358,  443,  687,  752, 1039, 1113, 1359, 1443, 2048+1692,
 193,  246,  424,  545,  564,  633,  828, 1047, 1323, 1324, 1400, 1532, 2048+1693,
   6,  380,  436,  467,  554,  611,  620,  621,  982, 1269, 1303, 1520, 2048+1694,
 313,  399,  656,  676,  695,  721,  762,  774,  851, 1310, 1325, 1545, 2048+1695,
  16,  497,  576,  577,  722,  753,  829,  905,  970, 1072, 1444, 1492, 2048+1696,
  69,  105,  301,  612,  634,  708, 1258, 1326, 1334, 1422, 1478, 1567, 2048+1697,
   7,  170,  280,  366,  498,  873,  917, 1080, 1201, 1213, 1278, 1378, 2048+1698,
 171,  457,  510,  534,  546,  688,  743,  786, 1061, 1081, 1114, 1546, 2048+1699,
 247,  400,  596,  641,  787, 1016, 1137, 1202, 1214, 1436, 1455, 1577, 2048+1700,
  60,  268,  314,  401,  478,  556,  642,  885,  950, 1238, 1311, 1558, 2048+1719,
  17,  147,  391,  444,  622,  744,  763,  831, 1026, 1246, 1521, 1522, 2048+1720,
 136,  204,  579,  635,  666,  754,  810,  818,  819, 1181, 1468, 1502, 2048+1721,
 161,  512,  598,  854,  875,  895,  920,  962,  972, 1049, 1510, 1523, 2048+1722,
  61,  107,  214,  696,  775,  776,  921,  951, 1027, 1104, 1169, 1270, 2048+1723,
  39,   93,  183,  269,  303,  499,  811,  832,  907, 1456, 1524, 1533, 2048+1724,
 205,  368,  479,  565,  697, 1073, 1115, 1279, 1401, 1413, 1479, 1578, 2048+1725,
 162,  369,  657,  709,  733,  745,  886,  941,  985, 1260, 1280, 1312, 2048+1726,
  51,   70,  194,  445,  599,  796,  841,  986, 1215, 1337, 1402, 1414, 2048+1727,
 173,  260,  468,  513,  600,  677,  756,  842, 1083, 1149, 1437, 1511, 2048+1746,
 137,  138,  215,  346,  590,  643,  820,  942,  963, 1029, 1225, 1445, 2048+1747,
  84,  118,  334,  402,  778,  833,  866,  952, 1008, 1018, 1019, 1379, 2048+1748,
 127,  139,  359,  711,  798, 1052, 1075, 1095, 1118, 1162, 1171, 1248, 2048+1749,
 261,  305,  414,  896,  973,  974, 1119, 1150, 1226, 1304, 1370, 1469, 2048+1750,
  71,  140,  148,  238,  293,  381,  469,  501,  698, 1009, 1030, 1106, 2048+1751,
  18,   28,   94,  195,  403,  567,  678,  764,  897, 1271, 1313, 1480, 2048+1752,
 360,  568,  855,  908,  932,  943, 1084, 1139, 1184, 1458, 1481, 1512, 2048+1753,
  19,   29,  250,  270,  392,  644,  799,  995, 1041, 1185, 1415, 1536, 2048+1754,
  52,  128,  371,  458,  667,  712,  800,  876,  954, 1042, 1282, 1349, 2048+1773,
  62,  335,  336,  415,  547,  789,  843, 1020, 1140, 1163, 1228, 1425, 2048+1774,
 283,  316,  536,  601,  976, 1031, 1064, 1151, 1206, 1217, 1218, 1579, 2048+1775,
 327,  337,  557,  910,  997, 1251, 1273, 1295, 1316, 1361, 1372, 1447, 2048+1776,
  85,  459,  503,  613, 1096, 1172, 1173, 1317, 1350, 1426, 1503, 1569, 2048+1777,
 271,  338,  347,  437,  492,  580,  668,  700,  898, 1207, 1229, 1306, 2048+1778,
  95,  216,  227,  294,  393,  602,  766,  877,  964, 1097, 1470, 1513, 2048+1779,
  73,   96,  129,  558,  767, 1053, 1107, 1130, 1141, 1283, 1339, 1382, 2048+1780,
  30,  151,  217,  228,  448,  470,  591,  844,  998, 1195, 1240, 1383, 2048+1781,

   8,   18, 2048+1440,
  19,   28, 2048+1441,
  29,   38, 2048+1442,
  39,   48, 2048+1443,
  49,   58, 2048+1444,
  59,   68, 2048+1445,
  69,   78, 2048+1446,
  79,   88, 2048+1447,
  89,   98, 2048+1448,
  99,  108, 2048+1449,
 109,  118, 2048+1450,
 119,  128, 2048+1451,
 129,  138, 2048+1452,
 139,  148, 2048+1453,
 149,  158, 2048+1454,
 159,  168, 2048+1455,
 169,  178, 2048+1456,
 179,  188, 2048+1457,
 189,  198, 2048+1458,
 199,  208, 2048+1459,
 209,  218, 2048+1460,
 219,  228, 2048+1461,
 229,  238, 2048+1462,
 239,  248, 2048+1463,
 249,  258, 2048+1464,
 259,  268, 2048+1465,
 269,  278, 2048+1466,
 279,  288, 2048+1467,
 289,  298, 2048+1468,
 299,  308, 2048+1469,
 309,  318, 2048+1470,
 319,  328, 2048+1471,
 329,  338, 2048+1472,
 339,  348, 2048+1473,
 349,  358, 2048+1474,
 359,  368, 2048+1475,
 369,  378, 2048+1476,
 379,  388, 2048+1477,
 389,  398, 2048+1478,
 399,  408, 2048+1479,
 409,  418, 2048+1480,
 419,  428, 2048+1481,
 429,  438, 2048+1482,
 439,  448, 2048+1483,
 449,  458, 2048+1484,
 459,  468, 2048+1485,
 469,  478, 2048+1486,
 479,  488, 2048+1487,
 489,  498, 2048+1488,
 499,  508, 2048+1489,
 509,  518, 2048+1490,
 519,  528, 2048+1491,
 529,  538, 2048+1492,
 539,  548, 2048+1493,
 549,  558, 2048+1494,
 559,  568, 2048+1495,
 569,  578, 2048+1496,
 579,  588, 2048+1497,
 589,  598, 2048+1498,
 599,  608, 2048+1499,
 609,  618, 2048+1500,
 619,  628, 2048+1501,
 629,  638, 2048+1502,
 639,  648, 2048+1503,
 649,  658, 2048+1504,
 659,  668, 2048+1505,
 669,  678, 2048+1506,
 679,  688, 2048+1507,
 689,  698, 2048+1508,
 699,  708, 2048+1509,
 709,  718, 2048+1510,
 719,  728, 2048+1511,
 729,  738, 2048+1512,
 739,  748, 2048+1513,
 749,  758, 2048+1514,
 759,  768, 2048+1515,
 769,  778, 2048+1516,
 779,  788, 2048+1517,
 789,  798, 2048+1518,
 799,  808, 2048+1519,
 809,  818, 2048+1520,
 819,  828, 2048+1521,
 829,  838, 2048+1522,
 839,  848, 2048+1523,
 849,  858, 2048+1524,
 859,  868, 2048+1525,
 869,  878, 2048+1526,
 879,  888, 2048+1527,
 889,  898, 2048+1528,
 899,  908, 2048+1529,
 909,  918, 2048+1530,
 919,  928, 2048+1531,
 929,  938, 2048+1532,
 939,  948, 2048+1533,
 949,  958, 2048+1534,
 959,  968, 2048+1535,
 969,  978, 2048+1536,
 979,  988, 2048+1537,
 989,  998, 2048+1538,
 999, 1008, 2048+1539,
1009, 1018, 2048+1540,
1019, 1028, 2048+1541,
1029, 1038, 2048+1542,
1039, 1048, 2048+1543,
1049, 1058, 2048+1544,
1059, 1068, 2048+1545,
1069, 1078, 2048+1546,
1079, 1088, 2048+1547,
1089, 1098, 2048+1548,
1099, 1108, 2048+1549,
1109, 1118, 2048+1550,
1119, 1128, 2048+1551,
1129, 1138, 2048+1552,
1139, 1148, 2048+1553,
1149, 1158, 2048+1554,
1159, 1168, 2048+1555,
1169, 1178, 2048+1556,
1179, 1188, 2048+1557,
1189, 1198, 2048+1558,
   9, 1199, 2048+1559,
  30,  491, 1021, 2048+1203,
  40, 1071, 1180, 2048+1204,
  51,  361,  800, 2048+1205,
  60,  241, 1100, 2048+1206,
  31,   71, 1022, 2048+1207,
  80,  111, 1160, 2048+1208,
  72,   91, 1120, 2048+1209,
 101,  430,  460, 2048+1210,
 112,  750, 1050, 2048+1211,
 120,  660,  850, 2048+1212,
  81,  131,  740, 2048+1213,
 140,  400,  630, 2048+1214,
   2,  160,  431, 2048+1215,
  11,  631, 1000, 2048+1216,
  22,  290, 1023, 2048+1217,
  32,  450,  980, 2048+1218,
  41,  520,  770, 2048+1219,
  52,  420, 1150, 2048+1220,
  61,  560, 1072, 2048+1221,
  73,  960, 1060, 2048+1222,
   3,   74,   82, 2048+1223,
  92,  801,  861, 2048+1224,
 102,  291,  480, 2048+1225,
 113,  830,  840, 2048+1226,
 121,  350,  881, 2048+1227,
  42,  132, 1110, 2048+1228,
 141,  492,  540, 2048+1229,
 180,  641, 1171, 2048+1233,
  24,  133,  191, 2048+1234,
 202,  511,  950, 2048+1235,
  53,  210,  392, 2048+1236,
 181,  221, 1172, 2048+1237,
 114,  230,  261, 2048+1238,
  75,  222,  243, 2048+1239,
 251,  580,  610, 2048+1240,
   4,  262,  900, 2048+1241,
 270,  811, 1001, 2048+1242,
 231,  281,  891, 2048+1243,
 292,  550,  780, 2048+1244,
 152,  310,  581, 2048+1245,
 162,  781, 1151, 2048+1246,
 172,  442, 1173, 2048+1247,
 182,  601, 1131, 2048+1248,
 192,  670,  920, 2048+1249,
 103,  203,  570, 2048+1250,
  25,  211,  710, 2048+1251,
  12,  223, 1111, 2048+1252,
 153,  224,  232, 2048+1253,
 244,  951, 1011, 2048+1254,
 252,  443,  632, 2048+1255,
 263,  981,  990, 2048+1256,
 271,  500, 1031, 2048+1257,
  62,  193,  282, 2048+1258,
 293,  642,  690, 2048+1259,
 123,  330,  792, 2048+1263,
 174,  283,  341, 2048+1264,
 353,  662, 1101, 2048+1265,
 204,  362,  543, 2048+1266,
 124,  331,  371, 2048+1267,
 264,  381,  411, 2048+1268,
 225,  372,  394, 2048+1269,
 402,  730,  762, 2048+1270,
 154,  412, 1051, 2048+1271,
 421,  962, 1152, 2048+1272,
 382,  433, 1041, 2048+1273,
 444,  701,  930, 2048+1274,
 302,  461,  731, 2048+1275,
 104,  312,  931, 2048+1276,
 125,  322,  592, 2048+1277,
  84,  332,  752, 2048+1278,
 342,  820, 1073, 2048+1279,
 253,  354,  720, 2048+1280,
 175,  363,  862, 2048+1281,
  63,  163,  373, 2048+1282,
 303,  374,  383, 2048+1283,
 395, 1102, 1162, 2048+1284,
 403,  593,  782, 2048+1285,
 413, 1132, 1140, 2048+1286,
 422,  650, 1182, 2048+1287,
 212,  343,  434, 2048+1288,
 445,  793,  841, 2048+1289,
 273,  481,  942, 2048+1293,
 324,  435,  494, 2048+1294,
  54,  503,  813, 2048+1295,
 355,  512,  693, 2048+1296,
 274,  482,  522, 2048+1297,
 414,  532,  562, 2048+1298,
 375,  523,  545, 2048+1299,
 552,  882,  913, 2048+1300,
   5,  304,  563, 2048+1301,
 105,  571, 1113, 2048+1302,
 533,  583, 1191, 2048+1303,
 594,  852, 1082, 2048+1304,
 453,  611,  883, 2048+1305,
 254,  463, 1083, 2048+1306,
 275,  473,  743, 2048+1307,
 234,  483,  902, 2048+1308,
  26,  495,  971, 2048+1309,
 404,  504,  871, 2048+1310,
 325,  513, 1012, 2048+1311,
 213,  313,  524, 2048+1312,
 454,  525,  534, 2048+1313,
  55,  116,  546, 2048+1314,
 553,  744,  932, 2048+1315,
  85,   93,  564, 2048+1316,
 135,  572,  802, 2048+1317,
 364,  496,  584, 2048+1318,
 595,  943,  991, 2048+1319,
 424,  633, 1092, 2048+1323,
 475,  585,  644, 2048+1324,
 205,  653,  964, 2048+1325,
 505,  663,  844, 2048+1326,
 425,  634,  672, 2048+1327,
 565,  682,  712, 2048+1328,
 526,  673,  695, 2048+1329,
 703, 1032, 1064, 2048+1330,
 155,  455,  713, 2048+1331,
  65,  255,  721, 2048+1332,
 143,  683,  733, 2048+1333,
  35,  745, 1003, 2048+1334,
 604,  763, 1033, 2048+1335,
  36,  405,  613, 2048+1336,
 426,  623,  894, 2048+1337,
 385,  635, 1053, 2048+1338,
 176,  645, 1122, 2048+1339,
 554,  654, 1025, 2048+1340,
 476,  664, 1163, 2048+1341,
 365,  464,  674, 2048+1342,
 605,  675,  684, 2048+1343,
 206,  266,  696, 2048+1344,
 704,  895, 1084, 2048+1345,
 235,  245,  714, 2048+1346,
 285,  722,  952, 2048+1347,
 514,  646,  734, 2048+1348,
 746, 1093, 1141, 2048+1349,
  45,  574,  783, 2048+1353,
 625,  735,  795, 2048+1354,
 356,  805, 1115, 2048+1355,
 655,  814,  994, 2048+1356,
 575,  784,  822, 2048+1357,
 715,  833,  864, 2048+1358,
 676,  823,  846, 2048+1359,
  16,  854, 1183, 2048+1360,
 305,  606,  865, 2048+1361,
 215,  406,  872, 2048+1362,
 295,  834,  885, 2048+1363,
 185,  896, 1154, 2048+1364,
 755,  914, 1184, 2048+1365,
 186,  555,  765, 2048+1366,
 576,  774, 1044, 2048+1367,
   7,  536,  785, 2048+1368,
  77,  326,  796, 2048+1369,
 705,  806, 1175, 2048+1370,
 117,  626,  815, 2048+1371,
 515,  614,  824, 2048+1372,
 756,  825,  835, 2048+1373,
 357,  416,  847, 2048+1374,
  37,  855, 1045, 2048+1375,
 386,  396,  866, 2048+1376,
 437,  873, 1103, 2048+1377,
 665,  797,  886, 2048+1378,
  46,   94,  897, 2048+1379,
 196,  724,  933, 2048+1383,
 776,  887,  945, 2048+1384,
  67,  506,  955, 2048+1385,
 807,  965, 1144, 2048+1386,
 725,  934,  973, 2048+1387,
 867,  984, 1014, 2048+1388,
 826,  974,  996, 2048+1389,
 136,  167, 1005, 2048+1390,
 456,  757, 1015, 2048+1391,
 367,  556, 1026, 2048+1392,
 447,  985, 1035, 2048+1393,
 107,  335, 1046, 2048+1394,
 137,  905, 1065, 2048+1395,
 336,  706,  916, 2048+1396,
 726,  924, 1194, 2048+1397,
 157,  686,  935, 2048+1398,
 227,  477,  946, 2048+1399,
 127,  856,  956, 2048+1400,
 267,  777,  966, 2048+1401,
 666,  766,  975, 2048+1402,
 906,  976,  986, 2048+1403,
 507,  567,  997, 2048+1404,
 187, 1006, 1195, 2048+1405,
 537,  547, 1016, 2048+1406,
  56,  587, 1027, 2048+1407,
 816,  947, 1036, 2048+1408,
 197,  246, 1047, 2048+1409,
 346,  875, 1085, 2048+1413,
 926, 1037, 1095, 2048+1414,
 217,  656, 1106, 2048+1415,
  97,  957, 1116, 2048+1416,
 876, 1086, 1124, 2048+1417,
1017, 1135, 1165, 2048+1418,
 977, 1125, 1146, 2048+1419,
 286,  317, 1156, 2048+1420,
 607,  907, 1166, 2048+1421,
 517,  707, 1176, 2048+1422,
 597, 1136, 1186, 2048+1423,
 257,  486, 1196, 2048+1424,
  17,  287, 1056, 2048+1425,
 487,  857, 1067, 2048+1426,
 146,  877, 1077, 2048+1427,
 307,  837, 1087, 2048+1428,
 377,  627, 1096, 2048+1429,
 277, 1007, 1107, 2048+1430,
 417,  927, 1117, 2048+1431,
 817,  917, 1126, 2048+1432,
1057, 1127, 1137, 2048+1433,
 657,  717, 1147, 2048+1434,
 147,  337, 1157, 2048+1435,
 687,  697, 1167, 2048+1436,
 207,  737, 1177, 2048+1437,
 967, 1097, 1187, 2048+1438,
 347,  397, 1197, 2048+1439,
   0,   90,  200,  440,  530,  600,  760,  810,  860,  910,  970, 1020, 1080, 2048+1200,
   1,   10,   20,  110,  130,  380,  470,  490,  761,  790,  870,  880, 1081, 2048+1201,
  21,   50,   70,  100,  190,  240,  360,  390,  441,  700,  890, 1070, 1130, 2048+1202,
  33,  150,  242,  351,  590,  680,  751,  911,  961, 1010, 1061, 1121, 1170, 2048+1230,
  34,  151,  161,  170,  260,  280,  531,  620,  640,  912,  940, 1024, 1030, 2048+1231,
  23,   83,  171,  201,  220,  250,  340,  391,  510,  541,  591,  851, 1040, 2048+1232,
  13,   76,  122,  183,  300,  393,  501,  741,  831,  901, 1062, 1112, 1161, 2048+1260,
 184,  301,  311,  320,  410,  432,  681,  771,  791, 1063, 1090, 1174, 1181, 2048+1261,
 173,  233,  321,  352,  370,  401,  493,  542,  661,  691,  742, 1002, 1190, 2048+1262,
  14,   64,  115,  164,  226,  272,  333,  451,  544,  651,  892,  982, 1052, 2048+1290,
  15,   43,  126,  134,  334,  452,  462,  471,  561,  582,  832,  921,  941, 2048+1291,
 142,  323,  384,  472,  502,  521,  551,  643,  692,  812,  842,  893, 1153, 2048+1292,
   6,  165,  214,  265,  314,  376,  423,  484,  602,  694,  803, 1042, 1133, 2048+1320,
 166,  194,  276,  284,  485,  603,  612,  621,  711,  732,  983, 1074, 1091, 2048+1321,
 106,  294,  474,  535,  622,  652,  671,  702,  794,  843,  963,  992, 1043, 2048+1322,
  86,  156,  315,  366,  415,  465,  527,  573,  636,  753,  845,  953, 1192, 2048+1350,
  27,   44,  316,  344,  427,  436,  637,  754,  764,  772,  863,  884, 1134, 2048+1351,
 256,  446,  624,  685,  773,  804,  821,  853,  944,  993, 1114, 1142, 1193, 2048+1352,
 144,  236,  306,  466,  516,  566,  615,  677,  723,  786,  903,  995, 1104, 2048+1380,
  87,  177,  195,  467,  497,  577,  586,  787,  904,  915,  922, 1013, 1034, 2048+1381,
  66,   95,  145,  407,  596,  775,  836,  923,  954,  972, 1004, 1094, 1143, 2048+1382,
  57,  296,  387,  457,  616,  667,  716,  767,  827,  874,  936, 1054, 1145, 2048+1410,
 237,  327,  345,  617,  647,  727,  736,  937, 1055, 1066, 1075, 1164, 1185, 2048+1411,
  47,   96,  216,  247,  297,  557,  747,  925,  987, 1076, 1105, 1123, 1155, 2048+1412,

   8,   20, 2048+1320,
  21,   31, 2048+1321,
  32,   40, 2048+1322,
  41,   50, 2048+1323,
  51,   63, 2048+1324,
  64,   74, 2048+1325,
  75,   86, 2048+1326,
  87,   97, 2048+1327,
  98,  107, 2048+1328,
 108,  118, 2048+1329,
 119,  130, 2048+1330,
 131,  140, 2048+1331,
 141,  152, 2048+1332,
 153,  163, 2048+1333,
 164,  172, 2048+1334,
 173,  182, 2048+1335,
 183,  195, 2048+1336,
 196,  206, 2048+1337,
 207,  218, 2048+1338,
 219,  229, 2048+1339,
 230,  239, 2048+1340,
 240,  250, 2048+1341,
 251,  262, 2048+1342,
 263,  272, 2048+1343,
 273,  284, 2048+1344,
 285,  295, 2048+1345,
 296,  304, 2048+1346,
 305,  314, 2048+1347,
 315,  327, 2048+1348,
 328,  338, 2048+1349,
 339,  350, 2048+1350,
 351,  361, 2048+1351,
 362,  371, 2048+1352,
 372,  382, 2048+1353,
 383,  394, 2048+1354,
 395,  404, 2048+1355,
 405,  416, 2048+1356,
 417,  427, 2048+1357,
 428,  436, 2048+1358,
 437,  446, 2048+1359,
 447,  459, 2048+1360,
 460,  470, 2048+1361,
 471,  482, 2048+1362,
 483,  493, 2048+1363,
 494,  503, 2048+1364,
 504,  514, 2048+1365,
 515,  526, 2048+1366,
 527,  536, 2048+1367,
 537,  548, 2048+1368,
 549,  559, 2048+1369,
 560,  568, 2048+1370,
 569,  578, 2048+1371,
 579,  591, 2048+1372,
 592,  602, 2048+1373,
 603,  614, 2048+1374,
 615,  625, 2048+1375,
 626,  635, 2048+1376,
 636,  646, 2048+1377,
 647,  658, 2048+1378,
 659,  668, 2048+1379,
 669,  680, 2048+1380,
 681,  691, 2048+1381,
 692,  700, 2048+1382,
 701,  710, 2048+1383,
 711,  723, 2048+1384,
 724,  734, 2048+1385,
 735,  746, 2048+1386,
 747,  757, 2048+1387,
 758,  767, 2048+1388,
 768,  778, 2048+1389,
 779,  790, 2048+1390,
 791,  800, 2048+1391,
 801,  812, 2048+1392,
 813,  823, 2048+1393,
 824,  832, 2048+1394,
 833,  842, 2048+1395,
 843,  855, 2048+1396,
 856,  866, 2048+1397,
 867,  878, 2048+1398,
 879,  889, 2048+1399,
 890,  899, 2048+1400,
 900,  910, 2048+1401,
 911,  922, 2048+1402,
 923,  932, 2048+1403,
 933,  944, 2048+1404,
 945,  955, 2048+1405,
 956,  964, 2048+1406,
 965,  974, 2048+1407,
 975,  987, 2048+1408,
 988,  998, 2048+1409,
 999, 1010, 2048+1410,
1011, 1021, 2048+1411,
1022, 1031, 2048+1412,
1032, 1042, 2048+1413,
1043, 1054, 2048+1414,
   9, 1055, 2048+1415,
  43,  252,  976, 2048+1057,
  52,  384, 1000, 2048+1058,
  65,  142,  495, 2048+1059,
  76,  946,  977, 2048+1060,
  10,   88,  484, 2048+1061,
  99,  593,  616, 2048+1062,
 109,  110,  154, 2048+1063,
 121,  265,  340, 2048+1064,
   0,  197,  604, 2048+1065,
  11,  297,  880, 2048+1066,
  22,  891,  924, 2048+1067,
  34,  396,  845, 2048+1068,
  44,  682,  978, 2048+1069,
  53,  505,  957, 2048+1070,
  66,  100,  881, 2048+1071,
  77,  506,  683, 2048+1072,
  89,  274,  605, 2048+1073,
 101,  306,  307, 2048+1074,
 111,  330,  385, 2048+1075,
 122,  143,  912, 2048+1076,
   1,   78,  882, 2048+1077,
  12,  352,  496, 2048+1078,
  23,  386,  449, 2048+1079,
  35,  406,  693, 2048+1080,
  13,   45,  208, 2048+1081,
  54,  286,  594, 2048+1082,
  67,  397,  507, 2048+1083,
  55,   79,  637, 2048+1084,
  90,  550,  627, 2048+1085,
 102,  429,  857, 2048+1086,
 112,  174,  438, 2048+1087,
 123,  266,  780, 2048+1088,
  56,  176,  387, 2048+1090,
  80,  184,  516, 2048+1091,
 198,  275,  628, 2048+1092,
  24,   57,  209, 2048+1093,
 144,  220,  617, 2048+1094,
 231,  725,  748, 2048+1095,
 241,  242,  287, 2048+1096,
 254,  399,  472, 2048+1097,
 132,  331,  736, 2048+1098,
 145,  430, 1012, 2048+1099,
   2,  155, 1023, 2048+1100,
 166,  528,  980, 2048+1101,
  58,  177,  815, 2048+1102,
  36,  185,  638, 2048+1103,
 199,  232, 1013, 2048+1104,
 210,  639,  816, 2048+1105,
 221,  407,  737, 2048+1106,
 233,  439,  440, 2048+1107,
 243,  462,  517, 2048+1108,
 255,  276, 1044, 2048+1109,
 133,  211, 1014, 2048+1110,
 146,  485,  629, 2048+1111,
 156,  518,  581, 2048+1112,
 167,  539,  825, 2048+1113,
 147,  178,  341, 2048+1114,
 186,  418,  726, 2048+1115,
 200,  529,  640, 2048+1116,
 187,  212,  769, 2048+1117,
 222,  684,  759, 2048+1118,
 234,  561,  989, 2048+1119,
 244,  308,  570, 2048+1120,
 256,  400,  913, 2048+1121,
 188,  310,  519, 2048+1123,
 213,  316,  648, 2048+1124,
 332,  408,  760, 2048+1125,
 157,  189,  342, 2048+1126,
 277,  353,  749, 2048+1127,
 363,  858,  883, 2048+1128,
 373,  374,  419, 2048+1129,
 389,  531,  606, 2048+1130,
 267,  463,  869, 2048+1131,
  91,  278,  562, 2048+1132,
 103,  134,  288, 2048+1133,
  60,  299,  660, 2048+1134,
 190,  311,  948, 2048+1135,
 168,  317,  770, 2048+1136,
  92,  333,  364, 2048+1137,
 343,  771,  949, 2048+1138,
 354,  540,  870, 2048+1139,
 365,  571,  572, 2048+1140,
 375,  596,  649, 2048+1141,
 124,  390,  409, 2048+1142,
  93,  268,  344, 2048+1143,
 279,  618,  761, 2048+1144,
 289,  650,  713, 2048+1145,
 300,  671,  958, 2048+1146,
 280,  312,  473, 2048+1147,
 318,  551,  859, 2048+1148,
 334,  661,  772, 2048+1149,
 319,  345,  901, 2048+1150,
 355,  817,  892, 2048+1151,
  68,  366,  694, 2048+1152,
 376,  441,  702, 2048+1153,
 391,  532, 1045, 2048+1154,
 320,  443,  651, 2048+1156,
 346,  450,  781, 2048+1157,
 464,  541,  893, 2048+1158,
 290,  321,  474, 2048+1159,
 410,  486,  884, 2048+1160,
 497,  990, 1015, 2048+1161,
 508,  509,  552, 2048+1162,
 521,  663,  738, 2048+1163,
 401,  597, 1002, 2048+1164,
 223,  411,  695, 2048+1165,
 235,  269,  420, 2048+1166,
 192,  432,  792, 2048+1167,
  26,  322,  444, 2048+1168,
 301,  451,  902, 2048+1169,
 224,  465,  498, 2048+1170,
  27,  475,  903, 2048+1171,
 487,  672, 1003, 2048+1172,
 499,  703,  704, 2048+1173,
 510,  728,  782, 2048+1174,
 257,  522,  542, 2048+1175,
 225,  402,  476, 2048+1176,
 412,  750,  894, 2048+1177,
 421,  783,  847, 2048+1178,
  37,  433,  804, 2048+1179,
 413,  445,  607, 2048+1180,
 452,  685,  991, 2048+1181,
 466,  793,  904, 2048+1182,
 453,  477, 1034, 2048+1183,
 488,  950, 1024, 2048+1184,
 201,  500,  826, 2048+1185,
 511,  573,  834, 2048+1186,
 125,  523,  664, 2048+1187,
 454,  575,  784, 2048+1189,
 478,  582,  914, 2048+1190,
 598,  673, 1025, 2048+1191,
 422,  455,  608, 2048+1192,
 543,  619, 1016, 2048+1193,
  69,   94,  630, 2048+1194,
 641,  642,  686, 2048+1195,
 653,  795,  871, 2048+1196,
  82,  533,  729, 2048+1197,
 356,  544,  827, 2048+1198,
 367,  403,  553, 2048+1199,
 324,  564,  925, 2048+1200,
 159,  456,  576, 2048+1201,
 434,  583, 1035, 2048+1202,
 357,  599,  631, 2048+1203,
 160,  609, 1036, 2048+1204,
  83,  620,  805, 2048+1205,
 632,  835,  836, 2048+1206,
 643,  861,  915, 2048+1207,
 392,  654,  674, 2048+1208,
 358,  534,  610, 2048+1209,
 545,  885, 1026, 2048+1210,
 554,  916,  982, 2048+1211,
 169,  565,  936, 2048+1212,
 546,  577,  739, 2048+1213,
  70,  584,  818, 2048+1214,
 600,  926, 1037, 2048+1215,
 114,  585,  611, 2048+1216,
  28,  104,  621, 2048+1217,
 335,  633,  959, 2048+1218,
 644,  705,  966, 2048+1219,
 258,  655,  796, 2048+1220,
 586,  707,  917, 2048+1222,
 612,  714, 1046, 2048+1223,
 105,  730,  806, 2048+1224,
 555,  587,  740, 2048+1225,
  95,  675,  751, 2048+1226,
 202,  226,  762, 2048+1227,
 773,  774,  819, 2048+1228,
 786,  928, 1004, 2048+1229,
 215,  665,  862, 2048+1230,
 489,  676,  960, 2048+1231,
 501,  535,  687, 2048+1232,
   3,  458,  697, 2048+1233,
 292,  588,  708, 2048+1234,
 115,  566,  715, 2048+1235,
 490,  731,  763, 2048+1236,
 116,  293,  741, 2048+1237,
 216,  752,  937, 2048+1238,
 764,  967,  968, 2048+1239,
 775,  993, 1047, 2048+1240,
 524,  787,  807, 2048+1241,
 491,  666,  742, 2048+1242,
 106,  677, 1017, 2048+1243,
  62,  688, 1048, 2048+1244,
  16,  302,  698, 2048+1245,
 678,  709,  872, 2048+1246,
 203,  716,  951, 2048+1247,
   4,  117,  732, 2048+1248,
 246,  717,  743, 2048+1249,
 161,  236,  753, 2048+1250,
  38,  467,  765, 2048+1251,
  46,  776,  837, 2048+1252,
 393,  788,  929, 2048+1253,
 718,  839, 1049, 2048+1255,
 126,  744,  848, 2048+1256,
 237,  863,  938, 2048+1257,
 689,  719,  873, 2048+1258,
 227,  808,  886, 2048+1259,
 336,  359,  895, 2048+1260,
 905,  906,  952, 2048+1261,
   6,   84,  919, 2048+1262,
 348,  797,  994, 2048+1263,
  39,  622,  809, 2048+1264,
 634,  667,  820, 2048+1265,
 135,  590,  829, 2048+1266,
 424,  720,  840, 2048+1267,
 247,  699,  849, 2048+1268,
 623,  864,  896, 2048+1269,
 248,  425,  874, 2048+1270,
  17,  349,  887, 2048+1271,
  47,   48,  897, 2048+1272,
  72,  127,  907, 2048+1273,
 656,  920,  939, 2048+1274,
 624,  798,  875, 2048+1275,
  96,  238,  810, 2048+1276,
 128,  194,  821, 2048+1277,
 150,  435,  830, 2048+1278,
 811,  841, 1005, 2048+1279,
  29,  337,  850, 2048+1280,
 136,  249,  865, 2048+1281,
 378,  851,  876, 2048+1282,
 294,  368,  888, 2048+1283,
 170,  601,  898, 2048+1284,
 179,  908,  969, 2048+1285,
   7,  525,  921, 2048+1286,
 129,  852,  971, 2048+1288,
 259,  877,  983, 2048+1289,
  18,  369,  995, 2048+1290,
 822,  853, 1006, 2048+1291,
 360,  940, 1018, 2048+1292,
 468,  492, 1027, 2048+1293,
  30, 1038, 1039, 2048+1294,
 138,  217, 1051, 2048+1295,
  73,  480,  930, 2048+1296,
 171,  754,  941, 2048+1297,
 766,  799,  953, 2048+1298,
 270,  722,  962, 2048+1299,
 557,  854,  972, 2048+1300,
 379,  831,  984, 2048+1301,
 755,  996, 1028, 2048+1302,
 380,  558, 1007, 2048+1303,
 151,  481, 1019, 2048+1304,
 180,  181, 1029, 2048+1305,
 205,  260, 1040, 2048+1306,
  19,  789, 1052, 2048+1307,
 756,  931, 1008, 2048+1308,
 228,  370,  942, 2048+1309,
 261,  326,  954, 2048+1310,
 283,  567,  963, 2048+1311,
  85,  943,  973, 2048+1312,
 162,  469,  985, 2048+1313,
 271,  381,  997, 2048+1314,
 513,  986, 1009, 2048+1315,
 426,  502, 1020, 2048+1316,
 303,  733, 1030, 2048+1317,
  49,  313, 1041, 2048+1318,
 139,  657, 1053, 2048+1319,
  33,   42,  120,  264,  329,  448,  538,  802,  814,  844,  868, 1033, 2048+1056,
 113,  165,  175,  253,  398,  461,  580,  670,  934,  947,  979, 1001, 2048+1089,
  14,   25,   59,   81,  245,  298,  309,  388,  530,  595,  712,  803, 2048+1122,
 148,  158,  191,  214,  377,  431,  442,  520,  662,  727,  846,  935, 2048+1155,
  15,  281,  291,  323,  347,  512,  563,  574,  652,  794,  860,  981, 2048+1188,
  61,  149,  414,  423,  457,  479,  645,  696,  706,  785,  927,  992, 2048+1221,
   5,   71,  193,  282,  547,  556,  589,  613,  777,  828,  838,  918, 2048+1254,
 137,  204,  325,  415,  679,  690,  721,  745,  909,  961,  970, 1050, 2048+1287,

  10,   21, 2048+1280,
  22,   34, 2048+1281,
  35,   46, 2048+1282,
  47,   58, 2048+1283,
  59,   71, 2048+1284,
  72,   84, 2048+1285,
  85,   97, 2048+1286,
  98,  110, 2048+1287,
 111,  123, 2048+1288,
 124,  135, 2048+1289,
 136,  146, 2048+1290,
 147,  159, 2048+1291,
 160,  171, 2048+1292,
 172,  183, 2048+1293,
 184,  196, 2048+1294,
 197,  209, 2048+1295,
 210,  222, 2048+1296,
 223,  235, 2048+1297,
 236,  248, 2048+1298,
 249,  260, 2048+1299,
 261,  271, 2048+1300,
 272,  284, 2048+1301,
 285,  296, 2048+1302,
 297,  308, 2048+1303,
 309,  321, 2048+1304,
 322,  334, 2048+1305,
 335,  347, 2048+1306,
 348,  360, 2048+1307,
 361,  373, 2048+1308,
 374,  385, 2048+1309,
 386,  396, 2048+1310,
 397,  409, 2048+1311,
 410,  421, 2048+1312,
 422,  433, 2048+1313,
 434,  446, 2048+1314,
 447,  459, 2048+1315,
 460,  472, 2048+1316,
 473,  485, 2048+1317,
 486,  498, 2048+1318,
 499,  510, 2048+1319,
 511,  521, 2048+1320,
 522,  534, 2048+1321,
 535,  546, 2048+1322,
 547,  558, 2048+1323,
 559,  571, 2048+1324,
 572,  584, 2048+1325,
 585,  597, 2048+1326,
 598,  610, 2048+1327,
 611,  623, 2048+1328,
 624,  635, 2048+1329,
 636,  646, 2048+1330,
 647,  659, 2048+1331,
 660,  671, 2048+1332,
 672,  683, 2048+1333,
 684,  696, 2048+1334,
 697,  709, 2048+1335,
 710,  722, 2048+1336,
 723,  735, 2048+1337,
 736,  748, 2048+1338,
 749,  760, 2048+1339,
 761,  771, 2048+1340,
 772,  784, 2048+1341,
 785,  796, 2048+1342,
 797,  808, 2048+1343,
 809,  821, 2048+1344,
 822,  834, 2048+1345,
 835,  847, 2048+1346,
 848,  860, 2048+1347,
 861,  873, 2048+1348,
 874,  885, 2048+1349,
 886,  896, 2048+1350,
 897,  909, 2048+1351,
 910,  921, 2048+1352,
 922,  933, 2048+1353,
 934,  946, 2048+1354,
 947,  959, 2048+1355,
 960,  972, 2048+1356,
 973,  985, 2048+1357,
 986,  998, 2048+1358,
  11,  999, 2048+1359,
  60,  198,  560, 2048+1000,
  73,  161,  298, 2048+1001,
  86,  125,  648, 2048+1002,
  87,   99,  737, 2048+1003,
 112,  649,  849, 2048+1004,
   0,  286,  336, 2048+1005,
  12,  685,  875, 2048+1006,
  23,  310,  923, 2048+1007,
  36,  536,  987, 2048+1008,
  48,  113,  773, 2048+1009,
  61,  375,  698, 2048+1010,
  74,  423,  573, 2048+1011,
  88,  850,  887, 2048+1012,
 100,  273,  851, 2048+1013,
 114,  762,  836, 2048+1014,
   1,  398,  961, 2048+1015,
   2,   13,  500, 2048+1016,
  24,  137,  852, 2048+1017,
  37,  810,  898, 2048+1018,
  49,  974,  988, 2048+1019,
  62,  287,  288, 2048+1020,
  75,  173,  948, 2048+1021,
  89,  512,  738, 2048+1022,
 101,  673,  711, 2048+1023,
 115,  185,  448, 2048+1024,
   3,   25,  798, 2048+1025,
  14,  513,  586, 2048+1026,
  26,  126,  763, 2048+1027,
  38,   39,  650, 2048+1028,
  50,  102,  739, 2048+1029,
  40,   63,  424, 2048+1030,
  76,  250,  811, 2048+1031,
  90,  612,  823, 2048+1032,
  77,  103,  837, 2048+1033,
 116,  311,  599, 2048+1034,
 186,  323,  686, 2048+1035,
 199,  289,  425, 2048+1036,
 211,  251,  774, 2048+1037,
 212,  224,  862, 2048+1038,
 237,  775,  975, 2048+1039,
 127,  411,  461, 2048+1040,
   4,  138,  812, 2048+1041,
  51,  148,  435, 2048+1042,
 117,  162,  661, 2048+1043,
 174,  238,  899, 2048+1044,
 187,  501,  824, 2048+1045,
 200,  548,  699, 2048+1046,
  15,  213,  976, 2048+1047,
 225,  399,  977, 2048+1048,
 239,  888,  962, 2048+1049,
  91,  128,  523, 2048+1050,
 129,  139,  625, 2048+1051,
 149,  262,  978, 2048+1052,
  27,  163,  935, 2048+1053,
 104,  118,  175, 2048+1054,
 188,  412,  413, 2048+1055,
  78,  201,  299, 2048+1056,
 214,  637,  863, 2048+1057,
 226,  799,  838, 2048+1058,
 240,  312,  574, 2048+1059,
 130,  150,  924, 2048+1060,
 140,  638,  712, 2048+1061,
 151,  252,  889, 2048+1062,
 164,  165,  776, 2048+1063,
 176,  227,  864, 2048+1064,
 166,  189,  549, 2048+1065,
 202,  376,  936, 2048+1066,
 215,  740,  949, 2048+1067,
 203,  228,  963, 2048+1068,
 241,  436,  724, 2048+1069,
 313,  449,  813, 2048+1070,
 324,  414,  550, 2048+1071,
 337,  377,  900, 2048+1072,
 338,  349,  989, 2048+1073,
 105,  362,  901, 2048+1074,
 253,  537,  587, 2048+1075,
 131,  263,  937, 2048+1076,
 177,  274,  561, 2048+1077,
 242,  290,  786, 2048+1078,
  28,  300,  363, 2048+1079,
 314,  626,  950, 2048+1080,
 325,  674,  825, 2048+1081,
 106,  141,  339, 2048+1082,
 107,  350,  524, 2048+1083,
  16,   92,  364, 2048+1084,
 216,  254,  651, 2048+1085,
 255,  264,  750, 2048+1086,
 108,  275,  387, 2048+1087,
  64,  152,  291, 2048+1088,
 229,  243,  301, 2048+1089,
 315,  538,  539, 2048+1090,
 204,  326,  426, 2048+1091,
 340,  764,  990, 2048+1092,
 351,  925,  964, 2048+1093,
 365,  437,  700, 2048+1094,
  52,  256,  276, 2048+1095,
 265,  765,  839, 2048+1096,
  17,  277,  378, 2048+1097,
 292,  293,  902, 2048+1098,
 302,  352,  991, 2048+1099,
 294,  316,  675, 2048+1100,
  65,  327,  502, 2048+1101,
  79,  341,  865, 2048+1102,
  93,  328,  353, 2048+1103,
 366,  562,  853, 2048+1104,
 438,  575,  938, 2048+1105,
 450,  540,  676, 2048+1106,
  29,  462,  503, 2048+1107,
 119,  463,  474, 2048+1108,
  30,  230,  487, 2048+1109,
 379,  662,  713, 2048+1110,
  66,  257,  388, 2048+1111,
 303,  400,  687, 2048+1112,
 367,  415,  911, 2048+1113,
 153,  427,  488, 2048+1114,
  80,  439,  751, 2048+1115,
 451,  800,  951, 2048+1116,
 231,  266,  464, 2048+1117,
 232,  475,  652, 2048+1118,
 142,  217,  489, 2048+1119,
 342,  380,  777, 2048+1120,
 381,  389,  876, 2048+1121,
 233,  401,  514, 2048+1122,
 190,  278,  416, 2048+1123,
 354,  368,  428, 2048+1124,
 440,  663,  664, 2048+1125,
 329,  452,  551, 2048+1126,
 120,  465,  890, 2048+1127,
  53,   94,  476, 2048+1128,
 490,  563,  826, 2048+1129,
 178,  382,  402, 2048+1130,
 390,  891,  965, 2048+1131,
 143,  403,  504, 2048+1132,
  31,  417,  418, 2048+1133,
 121,  429,  477, 2048+1134,
 419,  441,  801, 2048+1135,
 191,  453,  627, 2048+1136,
 205,  466,  992, 2048+1137,
 218,  454,  478, 2048+1138,
 491,  688,  979, 2048+1139,
  67,  564,  701, 2048+1140,
 576,  665,  802, 2048+1141,
 154,  588,  628, 2048+1142,
 244,  589,  600, 2048+1143,
 155,  355,  613, 2048+1144,
 505,  787,  840, 2048+1145,
 192,  383,  515, 2048+1146,
 430,  525,  814, 2048+1147,
  41,  492,  541, 2048+1148,
 279,  552,  614, 2048+1149,
 206,  565,  877, 2048+1150,
  81,  577,  926, 2048+1151,
 356,  391,  590, 2048+1152,
 357,  601,  778, 2048+1153,
 267,  343,  615, 2048+1154,
 467,  506,  903, 2048+1155,
   5,  507,  516, 2048+1156,
 358,  526,  639, 2048+1157,
 317,  404,  542, 2048+1158,
 479,  493,  553, 2048+1159,
 566,  788,  789, 2048+1160,
 455,  578,  677, 2048+1161,
  18,  245,  591, 2048+1162,
 179,  219,  602, 2048+1163,
 616,  689,  952, 2048+1164,
 304,  508,  527, 2048+1165,
  19,   95,  517, 2048+1166,
 268,  528,  629, 2048+1167,
 156,  543,  544, 2048+1168,
 246,  554,  603, 2048+1169,
 545,  567,  927, 2048+1170,
 318,  579,  752, 2048+1171,
 122,  330,  592, 2048+1172,
 344,  580,  604, 2048+1173,
 109,  617,  815, 2048+1174,
 193,  690,  827, 2048+1175,
 702,  790,  928, 2048+1176,
 280,  714,  753, 2048+1177,
 369,  715,  725, 2048+1178,
 281,  480,  741, 2048+1179,
 630,  912,  966, 2048+1180,
 319,  509,  640, 2048+1181,
 555,  653,  939, 2048+1182,
 167,  618,  666, 2048+1183,
 405,  678,  742, 2048+1184,
   6,  331,  691, 2048+1185,
  54,  207,  703, 2048+1186,
 481,  518,  716, 2048+1187,
 482,  726,  904, 2048+1188,
 392,  468,  743, 2048+1189,
  32,  593,  631, 2048+1190,
 132,  632,  641, 2048+1191,
 483,  654,  766, 2048+1192,
 442,  529,  667, 2048+1193,
 605,  619,  679, 2048+1194,
 692,  913,  914, 2048+1195,
 581,  704,  803, 2048+1196,
 144,  370,  717, 2048+1197,
 305,  345,  727, 2048+1198,
  82,  744,  816, 2048+1199,
 431,  633,  655, 2048+1200,
 145,  220,  642, 2048+1201,
 393,  656,  754, 2048+1202,
 282,  668,  669, 2048+1203,
 371,  680,  728, 2048+1204,
  55,  670,  693, 2048+1205,
 443,  705,  878, 2048+1206,
 247,  456,  718, 2048+1207,
 469,  706,  729, 2048+1208,
 234,  745,  940, 2048+1209,
 320,  817,  953, 2048+1210,
  56,  828,  915, 2048+1211,
 406,  841,  879, 2048+1212,
 494,  842,  854, 2048+1213,
 407,  606,  866, 2048+1214,
  42,   96,  755, 2048+1215,
 444,  634,  767, 2048+1216,
  68,  681,  779, 2048+1217,
 295,  746,  791, 2048+1218,
 530,  804,  867, 2048+1219,
 133,  457,  818, 2048+1220,
 180,  332,  829, 2048+1221,
 607,  643,  843, 2048+1222,
  33,  608,  855, 2048+1223,
 519,  594,  868, 2048+1224,
 157,  719,  756, 2048+1225,
 258,  757,  768, 2048+1226,
 609,  780,  892, 2048+1227,
 568,  657,  792, 2048+1228,
 730,  747,  805, 2048+1229,
  43,   44,  819, 2048+1230,
 707,  830,  929, 2048+1231,
 269,  495,  844, 2048+1232,
 432,  470,  856, 2048+1233,
 208,  869,  941, 2048+1234,
 556,  758,  781, 2048+1235,
 270,  346,  769, 2048+1236,
 520,  782,  880, 2048+1237,
 408,  793,  794, 2048+1238,
 496,  806,  857, 2048+1239,
 181,  795,  820, 2048+1240,
   7,  569,  831, 2048+1241,
 372,  582,  845, 2048+1242,
 595,  832,  858, 2048+1243,
  69,  359,  870, 2048+1244,
  83,  445,  942, 2048+1245,
  45,  182,  954, 2048+1246,
   8,  531,  967, 2048+1247,
 620,  968,  980, 2048+1248,
 532,  731,  993, 2048+1249,
 168,  221,  881, 2048+1250,
 570,  759,  893, 2048+1251,
 194,  807,  905, 2048+1252,
 420,  871,  916, 2048+1253,
 658,  930,  994, 2048+1254,
 259,  583,  943, 2048+1255,
 306,  458,  955, 2048+1256,
 732,  770,  969, 2048+1257,
 158,  733,  981, 2048+1258,
 644,  720,  995, 2048+1259,
 283,  846,  882, 2048+1260,
 384,  883,  894, 2048+1261,
  20,  734,  906, 2048+1262,
 694,  783,  917, 2048+1263,
 859,  872,  931, 2048+1264,
 169,  170,  944, 2048+1265,
  57,  833,  956, 2048+1266,
 394,  621,  970, 2048+1267,
 557,  596,  982, 2048+1268,
  70,  333,  996, 2048+1269,
 682,  884,  907, 2048+1270,
 395,  471,  895, 2048+1271,
   9,  645,  908, 2048+1272,
 533,  918,  919, 2048+1273,
 622,  932,  983, 2048+1274,
 307,  920,  945, 2048+1275,
 134,  695,  957, 2048+1276,
 497,  708,  971, 2048+1277,
 721,  958,  984, 2048+1278,
 195,  484,  997, 2048+1279,

  14,   30, 2048+1392,
  31,   46, 2048+1393,
  47,   62, 2048+1394,
  63,   81, 2048+1395,
  82,   99, 2048+1396,
 100,  118, 2048+1397,
 119,  135, 2048+1398,
 136,  151, 2048+1399,
 152,  167, 2048+1400,
 168,  183, 2048+1401,
 184,  199, 2048+1402,
 200,  218, 2048+1403,
 219,  236, 2048+1404,
 237,  255, 2048+1405,
 256,  272, 2048+1406,
 273,  288, 2048+1407,
 289,  304, 2048+1408,
 305,  320, 2048+1409,
 321,  336, 2048+1410,
 337,  355, 2048+1411,
 356,  373, 2048+1412,
 374,  392, 2048+1413,
 393,  409, 2048+1414,
 410,  425, 2048+1415,
 426,  441, 2048+1416,
 442,  457, 2048+1417,
 458,  473, 2048+1418,
 474,  492, 2048+1419,
 493,  510, 2048+1420,
 511,  529, 2048+1421,
 530,  546, 2048+1422,
 547,  562, 2048+1423,
 563,  578, 2048+1424,
 579,  594, 2048+1425,
 595,  610, 2048+1426,
 611,  629, 2048+1427,
 630,  647, 2048+1428,
 648,  666, 2048+1429,
 667,  683, 2048+1430,
 684,  699, 2048+1431,
 700,  715, 2048+1432,
 716,  731, 2048+1433,
 732,  747, 2048+1434,
 748,  766, 2048+1435,
 767,  784, 2048+1436,
 785,  803, 2048+1437,
 804,  820, 2048+1438,
 821,  836, 2048+1439,
 837,  852, 2048+1440,
 853,  868, 2048+1441,
 869,  884, 2048+1442,
 885,  903, 2048+1443,
 904,  921, 2048+1444,
 922,  940, 2048+1445,
 941,  957, 2048+1446,
 958,  973, 2048+1447,
 974,  989, 2048+1448,
 990, 1005, 2048+1449,
1006, 1021, 2048+1450,
1022, 1040, 2048+1451,
1041, 1058, 2048+1452,
1059, 1077, 2048+1453,
1078, 1094, 2048+1454,
  15, 1095, 2048+1455,
  64,  101,  257, 2048+1097,
  83,  137,  512, 2048+1098,
  32,  102,  169, 2048+1099,
 120,  338, 1042, 2048+1100,
   0,    1,  258, 2048+1101,
  16,  749,  786, 2048+1102,
  33,  564,  871, 2048+1103,
  49,  259,  822, 2048+1104,
  65,  306,  631, 2048+1105,
  66,   84,  650, 2048+1106,
 103,  768,  854, 2048+1107,
  50,  121,  290, 2048+1108,
   2,  494,  769, 2048+1109,
  17,  122,  702, 2048+1110,
  34,  274,  548, 2048+1111,
  51,  260,  991, 2048+1112,
  67,  339,  717, 2048+1113,
  85,  238,  459, 2048+1114,
 104,  838,  886, 2048+1115,
 123,  375,  733, 2048+1116,
   3,    4,  855, 2048+1117,
  18,  495,  770, 2048+1118,
  35,  703,  992, 2048+1119,
  52,  105,  154, 2048+1120,
  68,  261,  340, 2048+1121,
  86,  275,  872, 2048+1122,
 106,  873, 1060, 2048+1123,
 124,  612,  942, 2048+1124,
   5,   19,  496, 2048+1125,
  20,  596,  975, 2048+1126,
  36,  107,  443, 2048+1127,
  53,  108,  262, 2048+1128,
  69,   70,  170, 2048+1129,
  87,  412,  943, 2048+1130,
  88,  109,  597, 2048+1131,
 125,  341,  685, 2048+1132,
 204,  239,  394, 2048+1134,
 221,  276,  651, 2048+1135,
 171,  240,  307, 2048+1136,
  89,  263,  475, 2048+1137,
 138,  139,  395, 2048+1138,
 155,  887,  924, 2048+1139,
 172,  704, 1008, 2048+1140,
 186,  396,  959, 2048+1141,
 205,  444,  771, 2048+1142,
 206,  222,  788, 2048+1143,
 241,  906,  993, 2048+1144,
 187,  264,  427, 2048+1145,
 140,  632,  907, 2048+1146,
 156,  265,  840, 2048+1147,
 173,  413,  686, 2048+1148,
  37,  188,  397, 2048+1149,
 207,  476,  856, 2048+1150,
 223,  376,  598, 2048+1151,
 242,  976, 1023, 2048+1152,
 266,  513,  874, 2048+1153,
 141,  142,  994, 2048+1154,
 157,  633,  908, 2048+1155,
  38,  174,  841, 2048+1156,
 189,  243,  292, 2048+1157,
 208,  398,  477, 2048+1158,
 224,  414, 1009, 2048+1159,
 110,  244, 1010, 2048+1160,
 267,  750, 1079, 2048+1161,
 143,  158,  634, 2048+1162,
  21,  159,  734, 2048+1163,
 175,  245,  580, 2048+1164,
 190,  246,  399, 2048+1165,
 209,  210,  308, 2048+1166,
 225,  550, 1080, 2048+1167,
 226,  247,  735, 2048+1168,
 268,  478,  823, 2048+1169,
 345,  377,  531, 2048+1171,
 358,  415,  789, 2048+1172,
 309,  378,  445, 2048+1173,
 227,  400,  613, 2048+1174,
 277,  278,  532, 2048+1175,
 293, 1024, 1062, 2048+1176,
  55,  310,  842, 2048+1177,
   6,  323,  533, 2048+1178,
 346,  581,  909, 2048+1179,
 347,  359,  926, 2048+1180,
  39,  379, 1044, 2048+1181,
 324,  401,  565, 2048+1182,
 279,  772, 1045, 2048+1183,
 294,  402,  978, 2048+1184,
 311,  551,  824, 2048+1185,
 176,  325,  534, 2048+1186,
 348,  614,  995, 2048+1187,
 360,  514,  736, 2048+1188,
  22,   71,  380, 2048+1189,
 403,  652, 1011, 2048+1190,
  40,  280,  281, 2048+1191,
 295,  773, 1046, 2048+1192,
 177,  312,  979, 2048+1193,
 326,  381,  429, 2048+1194,
 349,  535,  615, 2048+1195,
  56,  361,  552, 2048+1196,
  57,  248,  382, 2048+1197,
 126,  404,  888, 2048+1198,
 282,  296,  774, 2048+1199,
 160,  297,  875, 2048+1200,
 313,  383,  718, 2048+1201,
 327,  384,  536, 2048+1202,
 350,  351,  446, 2048+1203,
 127,  362,  688, 2048+1204,
 363,  385,  876, 2048+1205,
 405,  616,  960, 2048+1206,
 482,  515,  668, 2048+1208,
 498,  553,  927, 2048+1209,
 447,  516,  582, 2048+1210,
 364,  537,  751, 2048+1211,
 416,  417,  669, 2048+1212,
  72,  112,  430, 2048+1213,
 192,  448,  980, 2048+1214,
 144,  461,  670, 2048+1215,
 483,  719, 1047, 2048+1216,
 484,  499, 1064, 2048+1217,
  91,  178,  517, 2048+1218,
 462,  538,  705, 2048+1219,
  92,  418,  910, 2048+1220,
  24,  431,  539, 2048+1221,
 449,  689,  961, 2048+1222,
 314,  463,  671, 2048+1223,
  41,  485,  752, 2048+1224,
 500,  653,  877, 2048+1225,
 161,  211,  518, 2048+1226,
  58,  540,  790, 2048+1227,
 179,  419,  420, 2048+1228,
  93,  432,  911, 2048+1229,
  25,  315,  450, 2048+1230,
 464,  519,  567, 2048+1231,
 486,  672,  753, 2048+1232,
 193,  501,  690, 2048+1233,
 194,  386,  520, 2048+1234,
 269,  541, 1025, 2048+1235,
 421,  433,  912, 2048+1236,
 298,  434, 1012, 2048+1237,
 451,  521,  857, 2048+1238,
 465,  522,  673, 2048+1239,
 487,  488,  583, 2048+1240,
 270,  502,  826, 2048+1241,
 503,  523, 1013, 2048+1242,
   7,  542,  754, 2048+1243,
 620,  654,  806, 2048+1245,
 636,  691, 1065, 2048+1246,
 584,  655,  720, 2048+1247,
 504,  674,  889, 2048+1248,
 554,  555,  807, 2048+1249,
 212,  250,  568, 2048+1250,
  26,  329,  585, 2048+1251,
 283,  600,  808, 2048+1252,
  94,  621,  858, 2048+1253,
 114,  622,  637, 2048+1254,
 229,  316,  656, 2048+1255,
 601,  675,  843, 2048+1256,
 230,  556, 1048, 2048+1257,
 163,  569,  676, 2048+1258,
   8,  586,  827, 2048+1259,
 452,  602,  809, 2048+1260,
 180,  623,  890, 2048+1261,
 638,  791, 1014, 2048+1262,
 299,  352,  657, 2048+1263,
 195,  677,  928, 2048+1264,
 317,  557,  558, 2048+1265,
 231,  570, 1049, 2048+1266,
 164,  453,  587, 2048+1267,
 603,  658,  707, 2048+1268,
 624,  810,  891, 2048+1269,
 330,  639,  828, 2048+1270,
 331,  524,  659, 2048+1271,
  73,  406,  678, 2048+1272,
 559,  571, 1050, 2048+1273,
  59,  435,  572, 2048+1274,
 588,  660,  996, 2048+1275,
 604,  661,  811, 2048+1276,
 625,  626,  721, 2048+1277,
 407,  640,  963, 2048+1278,
  60,  641,  662, 2048+1279,
 145,  679,  892, 2048+1280,
 758,  792,  945, 2048+1282,
 115,  776,  829, 2048+1283,
 722,  793,  859, 2048+1284,
 642,  812, 1026, 2048+1285,
 692,  693,  946, 2048+1286,
 353,  388,  708, 2048+1287,
 165,  467,  723, 2048+1288,
 422,  738,  947, 2048+1289,
 232,  759,  997, 2048+1290,
 252,  760,  777, 2048+1291,
 366,  454,  794, 2048+1292,
 739,  813,  981, 2048+1293,
  95,  367,  694, 2048+1294,
 301,  709,  814, 2048+1295,
 146,  724,  964, 2048+1296,
 589,  740,  948, 2048+1297,
 318,  761, 1027, 2048+1298,
  61,  778,  929, 2048+1299,
 436,  489,  795, 2048+1300,
 332,  815, 1066, 2048+1301,
 455,  695,  696, 2048+1302,
  96,  368,  710, 2048+1303,
 302,  590,  725, 2048+1304,
 741,  796,  845, 2048+1305,
 762,  949, 1028, 2048+1306,
 468,  779,  965, 2048+1307,
 469,  663,  797, 2048+1308,
 213,  543,  816, 2048+1309,
  97,  697,  711, 2048+1310,
 196,  573,  712, 2048+1311,
  42,  726,  798, 2048+1312,
 742,  799,  950, 2048+1313,
 763,  764,  860, 2048+1314,
  10,  544,  780, 2048+1315,
 197,  781,  800, 2048+1316,
 284,  817, 1029, 2048+1317,
 896,  930, 1082, 2048+1319,
 253,  914,  966, 2048+1320,
 861,  931,  998, 2048+1321,
  74,  782,  951, 2048+1322,
 830,  831, 1083, 2048+1323,
 490,  526,  846, 2048+1324,
 303,  606,  862, 2048+1325,
 560,  879, 1084, 2048+1326,
  43,  369,  897, 2048+1327,
 390,  898,  915, 2048+1328,
 506,  591,  932, 2048+1329,
  27,  880,  952, 2048+1330,
 233,  507,  832, 2048+1331,
 438,  847,  953, 2048+1332,
  11,  285,  863, 2048+1333,
 727,  881, 1085, 2048+1334,
  75,  456,  899, 2048+1335,
 198,  916, 1067, 2048+1336,
 574,  627,  933, 2048+1337,
 116,  470,  954, 2048+1338,
 592,  833,  834, 2048+1339,
 234,  508,  848, 2048+1340,
 439,  728,  864, 2048+1341,
 882,  934,  983, 2048+1342,
  76,  900, 1086, 2048+1343,
  12,  607,  917, 2048+1344,
 608,  801,  935, 2048+1345,
 354,  680,  955, 2048+1346,
 235,  835,  849, 2048+1347,
 333,  713,  850, 2048+1348,
 181,  865,  936, 2048+1349,
 883,  937, 1087, 2048+1350,
 901,  902,  999, 2048+1351,
 148,  681,  918, 2048+1352,
 334,  919,  938, 2048+1353,
  77,  423,  956, 2048+1354,
 129, 1033, 1068, 2048+1356,
  13,  391, 1052, 2048+1357,
  44, 1000, 1069, 2048+1358,
 214,  920, 1088, 2048+1359,
 130,  967,  968, 2048+1360,
 628,  665,  984, 2048+1361,
 440,  744, 1001, 2048+1362,
 131,  698, 1016, 2048+1363,
 182,  509, 1034, 2048+1364,
 528, 1035, 1053, 2048+1365,
 644,  729, 1070, 2048+1366,
 166, 1017, 1089, 2048+1367,
 370,  645,  969, 2048+1368,
 576,  985, 1090, 2048+1369,
 149,  424, 1002, 2048+1370,
 132,  866, 1018, 2048+1371,
 215,  593, 1036, 2048+1372,
 117,  335, 1054, 2048+1373,
 714,  765, 1071, 2048+1374,
 254,  609, 1091, 2048+1375,
 730,  970,  971, 2048+1376,
 371,  646,  986, 2048+1377,
 577,  867, 1003, 2048+1378,
  29, 1019, 1072, 2048+1379,
 133,  216, 1037, 2048+1380,
 150,  745, 1055, 2048+1381,
 746,  939, 1073, 2048+1382,
 491,  818, 1092, 2048+1383,
 372,  972,  987, 2048+1384,
 471,  851,  988, 2048+1385,
 319, 1004, 1074, 2048+1386,
 134, 1020, 1075, 2048+1387,
  45, 1038, 1039, 2048+1388,
 287,  819, 1056, 2048+1389,
 472, 1057, 1076, 2048+1390,
 217,  561, 1093, 2048+1391,
  48,  153,  201,  202,  203,  220,  411,  649,  701,  805,  870,  905,  923, 2048+1096,
 185,  291,  342,  343,  344,  357,  549,  787,  839,  944, 1007, 1043, 1061, 2048+1133,
  54,   90,  111,  322,  428,  479,  480,  481,  497,  687,  925,  977, 1081, 2048+1170,
  23,  128,  191,  228,  249,  460,  566,  617,  618,  619,  635,  825, 1063, 2048+1207,
 113,  162,  271,  328,  365,  387,  599,  706,  755,  756,  757,  775,  962, 2048+1244,
   9,  251,  300,  408,  466,  505,  525,  737,  844,  893,  894,  895,  913, 2048+1281,
 147,  389,  437,  545,  605,  643,  664,  878,  982, 1030, 1031, 1032, 1051, 2048+1318,
  28,   78,   79,   80,   98,  286,  527,  575,  682,  743,  783,  802, 1015, 2048+1355,

  25,   52, 2048+1400,
  53,   79, 2048+1401,
  80,  106, 2048+1402,
 107,  133, 2048+1403,
 134,  160, 2048+1404,
 161,  187, 2048+1405,
 188,  214, 2048+1406,
 215,  241, 2048+1407,
 242,  268, 2048+1408,
 269,  295, 2048+1409,
 296,  322, 2048+1410,
 323,  349, 2048+1411,
 350,  376, 2048+1412,
 377,  403, 2048+1413,
 404,  430, 2048+1414,
 431,  457, 2048+1415,
 458,  484, 2048+1416,
 485,  511, 2048+1417,
 512,  538, 2048+1418,
 539,  565, 2048+1419,
 566,  592, 2048+1420,
 593,  619, 2048+1421,
 620,  646, 2048+1422,
 647,  673, 2048+1423,
 674,  700, 2048+1424,
 701,  727, 2048+1425,
 728,  754, 2048+1426,
 755,  781, 2048+1427,
 782,  808, 2048+1428,
 809,  835, 2048+1429,
 836,  862, 2048+1430,
 863,  889, 2048+1431,
 890,  916, 2048+1432,
 917,  943, 2048+1433,
 944,  970, 2048+1434,
 971,  997, 2048+1435,
 998, 1024, 2048+1436,
1025, 1051, 2048+1437,
1052, 1078, 2048+1438,
  26, 1079, 2048+1439,
   1,  164,  486, 2048+1085,
  28,  379,  460, 2048+1086,
  56,  216,  837, 2048+1087,
  83,  271,  945, 2048+1088,
 109,  110,  324, 2048+1089,
   2,  217,  729, 2048+1090,
  29,  111,  756, 2048+1091,
  57,  165,  918, 2048+1092,
  84,  540,  946, 2048+1093,
 112,  432,  594, 2048+1094,
   3,  166,  568, 2048+1095,
  30,  461,  947, 2048+1096,
  58,   85,  462, 2048+1097,
  86,  351,  649, 2048+1098,
 113,  405,  783, 2048+1099,
   4,  244,  675, 2048+1100,
  31,  189,  838, 2048+1101,
  59,   60,   87, 2048+1102,
   5,   88, 1027, 2048+1103,
 114,  297, 1053, 2048+1104,
   6,   61,  487, 2048+1105,
  32,  406,  757, 2048+1106,
  62,  115,  569, 2048+1107,
  89,  650,  810, 2048+1108,
 116,  167,  865, 2048+1109,
   7,  758,  811, 2048+1110,
  33,  570,  651, 2048+1111,
  63,  117,  488, 2048+1112,
  90,  463,  866, 2048+1113,
 118,  948,  972, 2048+1114,
   8,    9,  839, 2048+1115,
  34,  218,  325, 2048+1116,
  64,  219,  245, 2048+1117,
  91,  702,  949, 2048+1118,
 119,  326,  652, 2048+1119,
 138,  300,  621, 2048+1125,
 169,  514,  596, 2048+1126,
 192,  352,  973, 2048+1127,
  10,  222,  408, 2048+1128,
 247,  248,  464, 2048+1129,
 139,  353,  867, 2048+1130,
 170,  249,  892, 2048+1131,
 193,  301, 1054, 2048+1132,
  11,  223,  676, 2048+1133,
 250,  571,  730, 2048+1134,
 140,  302,  704, 2048+1135,
  12,  171,  597, 2048+1136,
 194,  224,  598, 2048+1137,
 225,  489,  785, 2048+1138,
 251,  541,  919, 2048+1139,
 141,  381,  812, 2048+1140,
 172,  327,  974, 2048+1141,
 195,  196,  226, 2048+1142,
  93,  142,  227, 2048+1143,
 120,  252,  433, 2048+1144,
 143,  197,  622, 2048+1145,
 173,  542,  893, 2048+1146,
 198,  253,  705, 2048+1147,
 228,  786,  950, 2048+1148,
 254,  303, 1000, 2048+1149,
 144,  894,  951, 2048+1150,
 174,  706,  787, 2048+1151,
 199,  255,  623, 2048+1152,
 229,  599, 1001, 2048+1153,
  13,   35,  256, 2048+1154,
 145,  146,  975, 2048+1155,
 175,  354,  465, 2048+1156,
 200,  355,  382, 2048+1157,
  14,  230,  840, 2048+1158,
 257,  466,  788, 2048+1159,
 275,  436,  759, 2048+1165,
 305,  654,  732, 2048+1166,
  36,  330,  490, 2048+1167,
 147,  358,  544, 2048+1168,
 384,  385,  600, 2048+1169,
 276,  491, 1002, 2048+1170,
 306,  386, 1029, 2048+1171,
 121,  331,  437, 2048+1172,
 148,  359,  813, 2048+1173,
 387,  707,  868, 2048+1174,
 277,  438,  842, 2048+1175,
 149,  307,  733, 2048+1176,
 332,  360,  734, 2048+1177,
 361,  624,  921, 2048+1178,
 388,  677, 1055, 2048+1179,
 278,  516,  952, 2048+1180,
  37,  308,  467, 2048+1181,
 333,  334,  362, 2048+1182,
 232,  279,  363, 2048+1183,
 258,  389,  572, 2048+1184,
 280,  335,  760, 2048+1185,
 309,  678, 1030, 2048+1186,
 336,  390,  843, 2048+1187,
  15,  364,  922, 2048+1188,
  66,  391,  439, 2048+1189,
  16,  281, 1031, 2048+1190,
 310,  844,  923, 2048+1191,
 337,  392,  761, 2048+1192,
  67,  365,  735, 2048+1193,
 150,  176,  393, 2048+1194,
  38,  282,  283, 2048+1195,
 311,  492,  601, 2048+1196,
 338,  493,  517, 2048+1197,
 151,  366,  976, 2048+1198,
 394,  602,  924, 2048+1199,
 412,  575,  895, 2048+1205,
 441,  790,  870, 2048+1206,
 177,  470,  625, 2048+1207,
 284,  496,  680, 2048+1208,
 519,  520,  736, 2048+1209,
  68,  413,  626, 2048+1210,
  95,  442,  521, 2048+1211,
 259,  471,  576, 2048+1212,
 285,  497,  953, 2048+1213,
 522,  845, 1003, 2048+1214,
 414,  577,  978, 2048+1215,
 286,  443,  871, 2048+1216,
 472,  498,  872, 2048+1217,
 499,  762, 1057, 2048+1218,
 122,  523,  814, 2048+1219,
  17,  415,  656, 2048+1220,
 178,  444,  603, 2048+1221,
 473,  474,  500, 2048+1222,
 368,  416,  501, 2048+1223,
 395,  524,  708, 2048+1224,
 417,  475,  896, 2048+1225,
  96,  445,  815, 2048+1226,
 476,  525,  979, 2048+1227,
 152,  502, 1058, 2048+1228,
 202,  526,  578, 2048+1229,
  97,  153,  418, 2048+1230,
 446,  980, 1059, 2048+1231,
 477,  527,  897, 2048+1232,
 203,  503,  873, 2048+1233,
 287,  312,  528, 2048+1234,
 179,  419,  420, 2048+1235,
 447,  627,  737, 2048+1236,
 478,  628,  657, 2048+1237,
  39,  288,  504, 2048+1238,
 529,  738, 1060, 2048+1239,
 548,  711, 1032, 2048+1245,
 580,  926, 1005, 2048+1246,
 313,  606,  763, 2048+1247,
 421,  631,  817, 2048+1248,
 659,  660,  874, 2048+1249,
 204,  549,  764, 2048+1250,
 234,  581,  661, 2048+1251,
 396,  607,  712, 2048+1252,
  18,  422,  632, 2048+1253,
  69,  662,  981, 2048+1254,
  41,  550,  713, 2048+1255,
 423,  582, 1006, 2048+1256,
 608,  633, 1007, 2048+1257,
 124,  634,  898, 2048+1258,
 260,  663,  954, 2048+1259,
 154,  551,  792, 2048+1260,
 314,  583,  739, 2048+1261,
 609,  610,  635, 2048+1262,
 506,  552,  636, 2048+1263,
 530,  664,  846, 2048+1264,
 553,  611, 1033, 2048+1265,
 235,  584,  955, 2048+1266,
  42,  612,  665, 2048+1267,
 125,  289,  637, 2048+1268,
 340,  666,  714, 2048+1269,
 236,  290,  554, 2048+1270,
  43,  126,  585, 2048+1271,
 613,  667, 1034, 2048+1272,
 341,  638, 1008, 2048+1273,
 424,  448,  668, 2048+1274,
 315,  555,  556, 2048+1275,
 586,  765,  875, 2048+1276,
 614,  766,  793, 2048+1277,
 180,  425,  639, 2048+1278,
 127,  669,  876, 2048+1279,
  98,  684,  849, 2048+1285,
  71,  716, 1062, 2048+1286,
 449,  742,  899, 2048+1287,
 557,  769,  957, 2048+1288,
 795,  796, 1009, 2048+1289,
 342,  685,  900, 2048+1290,
 370,  717,  797, 2048+1291,
 531,  743,  850, 2048+1292,
 155,  558,  770, 2048+1293,
  44,  205,  798, 2048+1294,
 182,  686,  851, 2048+1295,
  72,  559,  718, 2048+1296,
  73,  744,  771, 2048+1297,
 262,  772, 1035, 2048+1298,
  19,  397,  799, 2048+1299,
 291,  687,  928, 2048+1300,
 450,  719,  877, 2048+1301,
 745,  746,  773, 2048+1302,
 641,  688,  774, 2048+1303,
 670,  800,  982, 2048+1304,
  99,  689,  747, 2048+1305,
  20,  371,  720, 2048+1306,
 183,  748,  801, 2048+1307,
 263,  426,  775, 2048+1308,
 480,  802,  852, 2048+1309,
 372,  427,  690, 2048+1310,
 184,  264,  721, 2048+1311,
 100,  749,  803, 2048+1312,
  74,  481,  776, 2048+1313,
 560,  587,  804, 2048+1314,
 451,  691,  692, 2048+1315,
 722,  901, 1010, 2048+1316,
 750,  902,  929, 2048+1317,
 316,  561,  777, 2048+1318,
 265,  805, 1011, 2048+1319,
 237,  821,  985, 2048+1325,
 129,  207,  854, 2048+1326,
 588,  880, 1036, 2048+1327,
  22,  693,  905, 2048+1328,
  75,  931,  932, 2048+1329,
 482,  822, 1037, 2048+1330,
 508,  855,  933, 2048+1331,
 671,  881,  986, 2048+1332,
 292,  694,  906, 2048+1333,
 185,  343,  934, 2048+1334,
 318,  823,  987, 2048+1335,
 208,  695,  856, 2048+1336,
 209,  882,  907, 2048+1337,
 101,  399,  908, 2048+1338,
 156,  532,  935, 2048+1339,
 428,  824, 1064, 2048+1340,
 589,  857, 1012, 2048+1341,
 883,  884,  909, 2048+1342,
 779,  825,  910, 2048+1343,
  45,  806,  936, 2048+1344,
 238,  826,  885, 2048+1345,
 157,  509,  858, 2048+1346,
 319,  886,  937, 2048+1347,
 400,  562,  911, 2048+1348,
 616,  938,  988, 2048+1349,
 510,  563,  827, 2048+1350,
 320,  401,  859, 2048+1351,
 239,  887,  939, 2048+1352,
 210,  617,  912, 2048+1353,
 696,  723,  940, 2048+1354,
 590,  828,  829, 2048+1355,
  76,  860, 1038, 2048+1356,
 888, 1039, 1065, 2048+1357,
 452,  697,  913, 2048+1358,
  77,  402,  941, 2048+1359,
  48,  373,  961, 2048+1365,
 267,  345,  990, 2048+1366,
 102,  724, 1015, 2048+1367,
 159,  830, 1042, 2048+1368,
 211, 1067, 1068, 2048+1369,
 103,  618,  962, 2048+1370,
 643,  991, 1069, 2048+1371,
  49,  807, 1016, 2048+1372,
 429,  831, 1043, 2048+1373,
 321,  483, 1070, 2048+1374,
  50,  454,  963, 2048+1375,
 346,  832,  992, 2048+1376,
 347, 1017, 1044, 2048+1377,
 240,  534, 1045, 2048+1378,
 293,  672, 1071, 2048+1379,
 131,  564,  964, 2048+1380,
  78,  725,  993, 2048+1381,
1018, 1019, 1046, 2048+1382,
 915,  965, 1047, 2048+1383,
 186,  942, 1072, 2048+1384,
 374,  966, 1020, 2048+1385,
 294,  644,  994, 2048+1386,
 455, 1021, 1073, 2048+1387,
 535,  698, 1048, 2048+1388,
  51,  752, 1074, 2048+1389,
 645,  699,  967, 2048+1390,
 456,  536,  995, 2048+1391,
 375, 1022, 1075, 2048+1392,
 348,  753, 1049, 2048+1393,
 833,  861, 1076, 2048+1394,
 726,  968,  969, 2048+1395,
 104,  212,  996, 2048+1396,
 105,  132, 1023, 2048+1397,
 591,  834, 1050, 2048+1398,
 213,  537, 1077, 2048+1399,
   0,  135,  864, 1026, 2048+1080,
  27,  270,  459,  891, 2048+1081,
  54,  243,  567,  648, 2048+1082,
  81,  162,  163,  378, 2048+1083,
  55,   82,  108,  136, 2048+1084,
  92,  137,  272,  999, 2048+1120,
 168,  407,  595, 1028, 2048+1121,
 190,  380,  703,  784, 2048+1122,
 220,  298,  299,  513, 2048+1123,
 191,  221,  246,  273, 2048+1124,
  65,  231,  274,  409, 2048+1160,
  94,  304,  543,  731, 2048+1161,
 328,  515,  841,  920, 2048+1162,
 356,  434,  435,  653, 2048+1163,
 329,  357,  383,  410, 2048+1164,
 201,  367,  411,  545, 2048+1200,
 233,  440,  679,  869, 2048+1201,
 468,  655,  977, 1056, 2048+1202,
 494,  573,  574,  789, 2048+1203,
 469,  495,  518,  546, 2048+1204,
 339,  505,  547,  681, 2048+1240,
 369,  579,  816, 1004, 2048+1241,
  40,  123,  604,  791, 2048+1242,
 629,  709,  710,  925, 2048+1243,
 605,  630,  658,  682, 2048+1244,
 479,  640,  683,  818, 2048+1280,
  70,  507,  715,  956, 2048+1281,
 181,  261,  740,  927, 2048+1282,
 767,  847,  848, 1061, 2048+1283,
 741,  768,  794,  819, 2048+1284,
 615,  778,  820,  958, 2048+1320,
  21,  206,  642,  853, 2048+1321,
 317,  398,  878, 1063, 2048+1322,
 128,  903,  983,  984, 2048+1323,
 879,  904,  930,  959, 2048+1324,
  23,  751,  914,  960, 2048+1360,
 158,  344,  780,  989, 2048+1361,
 130,  453,  533, 1013, 2048+1362,
  46,   47,  266, 1040, 2048+1363,
  24, 1014, 1041, 1066, 2048+1364);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , Do'length );
		end if;
	end process;
	
end Behavioral;