LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VNP_INPUT_FIFO is
	generic(
		z			: integer := 48;
		W			: integer := 8
	);
	Port (
		clk			: in  std_logic;
		
		WrEn		: in  std_logic;
		Din			: in  std_logic_vector(W*z-1 downto 0);
		
		RdEn		: in  std_logic;
		Dout		: out std_logic_vector(W*z-1 downto 0)
	);
end VNP_INPUT_FIFO;

architecture Behavioral of VNP_INPUT_FIFO is	
	type fifo_type is array (7 downto 0) of std_logic_vector(W*z-1 downto 0);
	signal fifo 		: fifo_type  := (others => (others => '0') );
	
	signal WrAddr		: std_logic_vector(2 downto 0) := (others => '0');
	signal RdAddr		: std_logic_vector(2 downto 0) := (others => '0');
begin
	process(clk)
	begin
		if rising_edge(clk) then
			if WrEn = '1' then
				WrAddr <= WrAddr + '1';
				fifo(conv_integer(WrAddr)) <= Din;
			end if;
			if RdEn = '1' then
				RdAddr <= RdAddr + '1';
			end if;
		end if;
	end process;
	Dout <= fifo(conv_integer(RdAddr));
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CNP_Input_Memory is
	Port (
		clk			: in  std_logic;
		
		RdAddr		: in  std_logic_vector(9 downto 0);
		Do			: out std_logic_vector(7 downto 0)
	);
end CNP_Input_Memory;

architecture Behavioral of CNP_Input_Memory is	
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 128*6-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
   0,  1,  2,  3,  4,  5+128
, 20, 21, 22, 23, 24, 25+128
, 26, 27, 28, 29, 30, 31+128
, 39, 40, 41, 42, 43, 44+128
, 45, 46, 47, 48, 49, 50+128
, 58, 59, 60, 61, 62, 63+128
, 64, 65, 66, 67, 68, 69+128
, 70, 71, 72, 73, 74, 75+128
,  6,  7,  8,  9, 10, 11, 12+128
, 13, 14, 15, 16, 17, 18, 19+128
, 32, 33, 34, 35, 36, 37, 38+128
, 51, 52, 53, 54, 55, 56, 57+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
,  0,  1,  2,  3,  4,  5,  6,  7,  8,  9+128
, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19+128
, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29+128
, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39+128
, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49+128
, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59+128
, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69+128
, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
,  0,  1,  2,  3,  4,  5,  6,  7,  8,  9+128
, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19+128
, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29+128
, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39+128
, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49+128
, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59+128
, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80+128
, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
,  0,  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13+128
, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27+128
, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41+128
, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70+128
, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84+128
, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
,  0,  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13+128
, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72+128
, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28+128
, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43+128
, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58+128
, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
,  0,  1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19+128
, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39+128
, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59+128
, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79+128
,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , 8 );
		end if;
	end process;
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CNP_Output_Memory is
	generic(
		z			: integer := 96
	);
	Port (
		clk			: in  std_logic;
		
		RdAddr		: in  std_logic_vector(9 downto 0);
		Do			: out std_logic_vector(13 downto 0)
	);
end CNP_Output_Memory;

architecture Behavioral of CNP_Output_Memory is	
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 128*6-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
(z-(94*z/96))*128+ 0, (z-(73*z/96))*128+ 1, (z-(55*z/96))*128+ 2, (z-(83*z/96))*128+ 3, (z-( 7*z/96))*128+ 4, (z-( 0*z/96))*128+ 5, 
(z-(61*z/96))*128+20, (z-(47*z/96))*128+21, (z-(65*z/96))*128+22, (z-(25*z/96))*128+23, (z-( 0*z/96))*128+24, (z-( 0*z/96))*128+25, 
(z-(39*z/96))*128+26, (z-(84*z/96))*128+27, (z-(41*z/96))*128+28, (z-(72*z/96))*128+29, (z-( 0*z/96))*128+30, (z-( 0*z/96))*128+31, 
(z-(95*z/96))*128+39, (z-(53*z/96))*128+40, (z-(14*z/96))*128+41, (z-(18*z/96))*128+42, (z-( 0*z/96))*128+43, (z-( 0*z/96))*128+44, 
(z-(11*z/96))*128+45, (z-(73*z/96))*128+46, (z-( 2*z/96))*128+47, (z-(47*z/96))*128+48, (z-( 0*z/96))*128+49, (z-( 0*z/96))*128+50, 
(z-(94*z/96))*128+58, (z-(59*z/96))*128+59, (z-(70*z/96))*128+60, (z-(72*z/96))*128+61, (z-( 0*z/96))*128+62, (z-( 0*z/96))*128+63, 
(z-( 7*z/96))*128+64, (z-(65*z/96))*128+65, (z-(39*z/96))*128+66, (z-(49*z/96))*128+67, (z-( 0*z/96))*128+68, (z-( 0*z/96))*128+69, 
(z-(43*z/96))*128+70, (z-(66*z/96))*128+71, (z-(41*z/96))*128+72, (z-(26*z/96))*128+73, (z-( 7*z/96))*128+74, (z-( 0*z/96))*128+75, 
(z-(27*z/96))*128+ 6, (z-(22*z/96))*128+ 7, (z-(79*z/96))*128+ 8, (z-( 9*z/96))*128+ 9, (z-(12*z/96))*128+10, (z-( 0*z/96))*128+11, (z-( 0*z/96))*128+12, 
(z-(24*z/96))*128+13, (z-(22*z/96))*128+14, (z-(81*z/96))*128+15, (z-(33*z/96))*128+16, (z-( 0*z/96))*128+17, (z-( 0*z/96))*128+18, (z-( 0*z/96))*128+19, 
(z-(46*z/96))*128+32, (z-(40*z/96))*128+33, (z-(82*z/96))*128+34, (z-(79*z/96))*128+35, (z-( 0*z/96))*128+36, (z-( 0*z/96))*128+37, (z-( 0*z/96))*128+38, 
(z-(12*z/96))*128+51, (z-(83*z/96))*128+52, (z-(24*z/96))*128+53, (z-(43*z/96))*128+54, (z-(51*z/96))*128+55, (z-( 0*z/96))*128+56, (z-( 0*z/96))*128+57, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
(z-( 3 mod z))*128+ 0, (z-( 0 mod z))*128+ 1, (z-( 2 mod z))*128+ 2, (z-( 0 mod z))*128+ 3, (z-( 3 mod z))*128+ 4, (z-( 7 mod z))*128+ 5, (z-( 1 mod z))*128+ 6, (z-( 1 mod z))*128+ 7, (z-( 1 mod z))*128+ 8, (z-( 0 mod z))*128+ 9, 
(z-( 1 mod z))*128+10, (z-(36 mod z))*128+11, (z-(34 mod z))*128+12, (z-(10 mod z))*128+13, (z-(18 mod z))*128+14, (z-( 2 mod z))*128+15, (z-( 3 mod z))*128+16, (z-( 0 mod z))*128+17, (z-( 0 mod z))*128+18, (z-( 0 mod z))*128+19, 
(z-(12 mod z))*128+20, (z-( 2 mod z))*128+21, (z-(15 mod z))*128+22, (z-(40 mod z))*128+23, (z-( 3 mod z))*128+24, (z-(15 mod z))*128+25, (z-( 2 mod z))*128+26, (z-(13 mod z))*128+27, (z-( 0 mod z))*128+28, (z-( 0 mod z))*128+29, 
(z-(19 mod z))*128+30, (z-(24 mod z))*128+31, (z-( 3 mod z))*128+32, (z-( 0 mod z))*128+33, (z-( 6 mod z))*128+34, (z-(17 mod z))*128+35, (z-( 8 mod z))*128+36, (z-(39 mod z))*128+37, (z-( 0 mod z))*128+38, (z-( 0 mod z))*128+39, 
(z-(20 mod z))*128+40, (z-( 6 mod z))*128+41, (z-(10 mod z))*128+42, (z-(29 mod z))*128+43, (z-(28 mod z))*128+44, (z-(14 mod z))*128+45, (z-(38 mod z))*128+46, (z-( 0 mod z))*128+47, (z-( 0 mod z))*128+48, (z-( 0 mod z))*128+49, 
(z-(10 mod z))*128+50, (z-(28 mod z))*128+51, (z-(20 mod z))*128+52, (z-( 8 mod z))*128+53, (z-(36 mod z))*128+54, (z-( 9 mod z))*128+55, (z-(21 mod z))*128+56, (z-(45 mod z))*128+57, (z-( 0 mod z))*128+58, (z-( 0 mod z))*128+59, 
(z-(35 mod z))*128+60, (z-(25 mod z))*128+61, (z-(37 mod z))*128+62, (z-(21 mod z))*128+63, (z-( 5 mod z))*128+64, (z-( 0 mod z))*128+65, (z-( 4 mod z))*128+66, (z-(20 mod z))*128+67, (z-( 0 mod z))*128+68, (z-( 0 mod z))*128+69, 
(z-( 6 mod z))*128+70, (z-( 6 mod z))*128+71, (z-( 4 mod z))*128+72, (z-(14 mod z))*128+73, (z-(30 mod z))*128+74, (z-( 3 mod z))*128+75, (z-(36 mod z))*128+76, (z-(14 mod z))*128+77, (z-( 1 mod z))*128+78, (z-( 0 mod z))*128+79, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
(z-( 2*z/96))*128+ 0, (z-(19*z/96))*128+ 1, (z-(47*z/96))*128+ 2, (z-(48*z/96))*128+ 3, (z-(36*z/96))*128+ 4, (z-(82*z/96))*128+ 5, (z-(47*z/96))*128+ 6, (z-(15*z/96))*128+ 7, (z-(95*z/96))*128+ 8, (z-( 0*z/96))*128+ 9, 
(z-(69*z/96))*128+10, (z-(88*z/96))*128+11, (z-(33*z/96))*128+12, (z-( 3*z/96))*128+13, (z-(16*z/96))*128+14, (z-(37*z/96))*128+15, (z-(40*z/96))*128+16, (z-(48*z/96))*128+17, (z-( 0*z/96))*128+18, (z-( 0*z/96))*128+19, 
(z-(10*z/96))*128+20, (z-(86*z/96))*128+21, (z-(62*z/96))*128+22, (z-(28*z/96))*128+23, (z-(85*z/96))*128+24, (z-(16*z/96))*128+25, (z-(34*z/96))*128+26, (z-(73*z/96))*128+27, (z-( 0*z/96))*128+28, (z-( 0*z/96))*128+29, 
(z-(28*z/96))*128+30, (z-(32*z/96))*128+31, (z-(81*z/96))*128+32, (z-(27*z/96))*128+33, (z-(88*z/96))*128+34, (z-( 5*z/96))*128+35, (z-(56*z/96))*128+36, (z-(37*z/96))*128+37, (z-( 0*z/96))*128+38, (z-( 0*z/96))*128+39, 
(z-(23*z/96))*128+40, (z-(29*z/96))*128+41, (z-(15*z/96))*128+42, (z-(30*z/96))*128+43, (z-(66*z/96))*128+44, (z-(24*z/96))*128+45, (z-(50*z/96))*128+46, (z-(62*z/96))*128+47, (z-( 0*z/96))*128+48, (z-( 0*z/96))*128+49, 
(z-(30*z/96))*128+50, (z-(65*z/96))*128+51, (z-(54*z/96))*128+52, (z-(14*z/96))*128+53, (z-( 0*z/96))*128+54, (z-(30*z/96))*128+55, (z-(74*z/96))*128+56, (z-( 0*z/96))*128+57, (z-( 0*z/96))*128+58, (z-( 0*z/96))*128+59, 
(z-( 0*z/96))*128+71, (z-(47*z/96))*128+72, (z-(13*z/96))*128+73, (z-(61*z/96))*128+74, (z-(84*z/96))*128+75, (z-(55*z/96))*128+76, (z-(78*z/96))*128+77, (z-(41*z/96))*128+78, (z-(95*z/96))*128+79, (z-( 0*z/96))*128+80, 
(z-(32*z/96))*128+60, (z-( 0*z/96))*128+61, (z-(15*z/96))*128+62, (z-(56*z/96))*128+63, (z-(85*z/96))*128+64, (z-( 5*z/96))*128+65, (z-( 6*z/96))*128+66, (z-(52*z/96))*128+67, (z-( 0*z/96))*128+68, (z-( 0*z/96))*128+69, (z-( 0*z/96))*128+70, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
(z-( 6*z/96))*128+ 0, (z-(38*z/96))*128+ 1, (z-( 3*z/96))*128+ 2, (z-(93*z/96))*128+ 3, (z-(30*z/96))*128+ 4, (z-(70*z/96))*128+ 5, (z-(86*z/96))*128+ 6, (z-(37*z/96))*128+ 7, (z-(38*z/96))*128+ 8, (z-( 4*z/96))*128+ 9, (z-(11*z/96))*128+10, (z-(46*z/96))*128+11, (z-(48*z/96))*128+12, (z-( 0*z/96))*128+13, 
(z-(62*z/96))*128+14, (z-(94*z/96))*128+15, (z-(19*z/96))*128+16, (z-(84*z/96))*128+17, (z-(92*z/96))*128+18, (z-(78*z/96))*128+19, (z-(15*z/96))*128+20, (z-(92*z/96))*128+21, (z-(45*z/96))*128+22, (z-(24*z/96))*128+23, (z-(32*z/96))*128+24, (z-(30*z/96))*128+25, (z-( 0*z/96))*128+26, (z-( 0*z/96))*128+27, 
(z-(71*z/96))*128+28, (z-(55*z/96))*128+29, (z-(12*z/96))*128+30, (z-(66*z/96))*128+31, (z-(45*z/96))*128+32, (z-(79*z/96))*128+33, (z-(78*z/96))*128+34, (z-(10*z/96))*128+35, (z-(22*z/96))*128+36, (z-(55*z/96))*128+37, (z-(70*z/96))*128+38, (z-(82*z/96))*128+39, (z-( 0*z/96))*128+40, (z-( 0*z/96))*128+41, 
(z-(32*z/96))*128+57, (z-(52*z/96))*128+58, (z-(55*z/96))*128+59, (z-(80*z/96))*128+60, (z-(95*z/96))*128+61, (z-(22*z/96))*128+62, (z-( 6*z/96))*128+63, (z-(51*z/96))*128+64, (z-(24*z/96))*128+65, (z-(90*z/96))*128+66, (z-(44*z/96))*128+67, (z-(20*z/96))*128+68, (z-( 0*z/96))*128+69, (z-( 0*z/96))*128+70, 
(z-(63*z/96))*128+71, (z-(31*z/96))*128+72, (z-(88*z/96))*128+73, (z-(20*z/96))*128+74, (z-( 6*z/96))*128+75, (z-(40*z/96))*128+76, (z-(56*z/96))*128+77, (z-(16*z/96))*128+78, (z-(71*z/96))*128+79, (z-(53*z/96))*128+80, (z-(27*z/96))*128+81, (z-(26*z/96))*128+82, (z-(48*z/96))*128+83, (z-( 0*z/96))*128+84, 
(z-(38*z/96))*128+42, (z-(61*z/96))*128+43, (z-(66*z/96))*128+44, (z-( 9*z/96))*128+45, (z-(73*z/96))*128+46, (z-(47*z/96))*128+47, (z-(64*z/96))*128+48, (z-(39*z/96))*128+49, (z-(61*z/96))*128+50, (z-(43*z/96))*128+51, (z-(95*z/96))*128+52, (z-(32*z/96))*128+53, (z-( 0*z/96))*128+54, (z-( 0*z/96))*128+55, (z-( 0*z/96))*128+56, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
(z-(81*z/96))*128+ 0, (z-(28*z/96))*128+ 1, (z-(14*z/96))*128+ 2, (z-(25*z/96))*128+ 3, (z-(17*z/96))*128+ 4, (z-(85*z/96))*128+ 5, (z-(29*z/96))*128+ 6, (z-(52*z/96))*128+ 7, (z-(78*z/96))*128+ 8, (z-(95*z/96))*128+ 9, (z-(22*z/96))*128+10, (z-(92*z/96))*128+11, (z-( 0*z/96))*128+12, (z-( 0*z/96))*128+13, 
(z-(53*z/96))*128+59, (z-(60*z/96))*128+60, (z-(80*z/96))*128+61, (z-(26*z/96))*128+62, (z-(75*z/96))*128+63, (z-(86*z/96))*128+64, (z-(77*z/96))*128+65, (z-( 1*z/96))*128+66, (z-( 3*z/96))*128+67, (z-(72*z/96))*128+68, (z-(60*z/96))*128+69, (z-(25*z/96))*128+70, (z-( 0*z/96))*128+71, (z-( 0*z/96))*128+72, 
(z-(42*z/96))*128+14, (z-(14*z/96))*128+15, (z-(68*z/96))*128+16, (z-(32*z/96))*128+17, (z-(70*z/96))*128+18, (z-(43*z/96))*128+19, (z-(11*z/96))*128+20, (z-(36*z/96))*128+21, (z-(40*z/96))*128+22, (z-(33*z/96))*128+23, (z-(57*z/96))*128+24, (z-(38*z/96))*128+25, (z-(24*z/96))*128+26, (z-( 0*z/96))*128+27, (z-( 0*z/96))*128+28, 
(z-(20*z/96))*128+29, (z-(63*z/96))*128+30, (z-(39*z/96))*128+31, (z-(70*z/96))*128+32, (z-(67*z/96))*128+33, (z-(38*z/96))*128+34, (z-( 4*z/96))*128+35, (z-(72*z/96))*128+36, (z-(47*z/96))*128+37, (z-(29*z/96))*128+38, (z-(60*z/96))*128+39, (z-( 5*z/96))*128+40, (z-(80*z/96))*128+41, (z-( 0*z/96))*128+42, (z-( 0*z/96))*128+43, 
(z-(64*z/96))*128+44, (z-( 2*z/96))*128+45, (z-(63*z/96))*128+46, (z-( 3*z/96))*128+47, (z-(51*z/96))*128+48, (z-(81*z/96))*128+49, (z-(15*z/96))*128+50, (z-(94*z/96))*128+51, (z-( 9*z/96))*128+52, (z-(85*z/96))*128+53, (z-(36*z/96))*128+54, (z-(14*z/96))*128+55, (z-(19*z/96))*128+56, (z-( 0*z/96))*128+57, (z-( 0*z/96))*128+58, 
(z-(77*z/96))*128+73, (z-(15*z/96))*128+74, (z-(28*z/96))*128+75, (z-(35*z/96))*128+76, (z-(72*z/96))*128+77, (z-(30*z/96))*128+78, (z-(68*z/96))*128+79, (z-(85*z/96))*128+80, (z-(84*z/96))*128+81, (z-(26*z/96))*128+82, (z-(64*z/96))*128+83, (z-(11*z/96))*128+84, (z-(89*z/96))*128+85, (z-( 0*z/96))*128+86, (z-( 0*z/96))*128+87, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
(z-( 1*z/96))*128+ 0, (z-(25*z/96))*128+ 1, (z-(55*z/96))*128+ 2, (z-(47*z/96))*128+ 3, (z-( 4*z/96))*128+ 4, (z-(91*z/96))*128+ 5, (z-(84*z/96))*128+ 6, (z-( 8*z/96))*128+ 7, (z-(86*z/96))*128+ 8, (z-(52*z/96))*128+ 9, (z-(82*z/96))*128+10, (z-(33*z/96))*128+11, (z-( 5*z/96))*128+12, (z-( 0*z/96))*128+13, (z-(36*z/96))*128+14, (z-(20*z/96))*128+15, (z-( 4*z/96))*128+16, (z-(77*z/96))*128+17, (z-(80*z/96))*128+18, (z-( 0*z/96))*128+19, 
(z-( 6*z/96))*128+20, (z-(36*z/96))*128+21, (z-(40*z/96))*128+22, (z-(47*z/96))*128+23, (z-(12*z/96))*128+24, (z-(79*z/96))*128+25, (z-(47*z/96))*128+26, (z-(41*z/96))*128+27, (z-(21*z/96))*128+28, (z-(12*z/96))*128+29, (z-(71*z/96))*128+30, (z-(14*z/96))*128+31, (z-(72*z/96))*128+32, (z-( 0*z/96))*128+33, (z-(44*z/96))*128+34, (z-(49*z/96))*128+35, (z-( 0*z/96))*128+36, (z-( 0*z/96))*128+37, (z-( 0*z/96))*128+38, (z-( 0*z/96))*128+39, 
(z-(51*z/96))*128+40, (z-(81*z/96))*128+41, (z-(83*z/96))*128+42, (z-( 4*z/96))*128+43, (z-(67*z/96))*128+44, (z-(21*z/96))*128+45, (z-(31*z/96))*128+46, (z-(24*z/96))*128+47, (z-(91*z/96))*128+48, (z-(61*z/96))*128+49, (z-(81*z/96))*128+50, (z-( 9*z/96))*128+51, (z-(86*z/96))*128+52, (z-(78*z/96))*128+53, (z-(60*z/96))*128+54, (z-(88*z/96))*128+55, (z-(67*z/96))*128+56, (z-(15*z/96))*128+57, (z-( 0*z/96))*128+58, (z-( 0*z/96))*128+59, 
(z-(50*z/96))*128+60, (z-(50*z/96))*128+61, (z-(15*z/96))*128+62, (z-(36*z/96))*128+63, (z-(13*z/96))*128+64, (z-(10*z/96))*128+65, (z-(11*z/96))*128+66, (z-(20*z/96))*128+67, (z-(53*z/96))*128+68, (z-(90*z/96))*128+69, (z-(29*z/96))*128+70, (z-(92*z/96))*128+71, (z-(57*z/96))*128+72, (z-(30*z/96))*128+73, (z-(84*z/96))*128+74, (z-(92*z/96))*128+75, (z-(11*z/96))*128+76, (z-(66*z/96))*128+77, (z-(80*z/96))*128+78, (z-( 0*z/96))*128+79, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)), 14);
		end if;
	end process;
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VNP_Input_Memory is
	Port (
		clk			: in  std_logic;
		
		RdAddr		: in  std_logic_vector(9 downto 0);
		Do			: out std_logic_vector(7 downto 0)
	);
end VNP_Input_Memory;

architecture Behavioral of VNP_Input_Memory is	
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 128*6-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
 5, 11, 117+128, 
12, 18, 118+128, 
19, 24, 119+128, 
25, 30, 120+128, 
31, 37, 121+128, 
38, 43, 122+128, 
44, 49, 123+128, 
50, 56, 124+128, 
57, 62, 125+128, 
63, 68, 126+128, 
69, 75, 127+128, 
20, 51, 70, 104+128, 
 0,  6, 45, 105+128, 
13, 40, 65, 107+128, 
14, 32, 52, 108+128, 
 8, 27, 47, 110+128, 
 2, 22, 66, 112+128, 
29, 42, 60, 114+128, 
 4, 36, 74, 116+128, 
 1, 21, 26, 39, 46, 64, 106+128, 
 7, 15, 33, 53, 58, 71, 109+128, 
 9, 16, 34, 54, 59, 72, 111+128, 
 3, 23, 28, 41, 48, 67, 113+128, 
10, 17, 35, 55, 61, 73, 115+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
 9, 18, 121+128, 
19, 28, 122+128, 
29, 38, 123+128, 
39, 48, 124+128, 
49, 58, 125+128, 
59, 68, 126+128, 
69, 79, 127+128, 
 0, 40, 60, 104+128, 
 1, 61, 70, 105+128, 
21, 31, 62, 107+128, 
 2, 11, 51, 108+128, 
33, 43, 72, 110+128, 
 4, 12, 23, 111+128, 
24, 44, 74, 113+128, 
 6, 35, 54, 114+128, 
15, 55, 76, 116+128, 
26, 46, 66, 117+128, 
17, 37, 57, 119+128, 
 8, 47, 78, 120+128, 
10, 20, 30, 41, 50, 71, 106+128, 
 3, 22, 32, 42, 52, 63, 109+128, 
 5, 13, 34, 53, 64, 73, 112+128, 
 7, 14, 25, 45, 65, 75, 115+128, 
16, 27, 36, 56, 67, 77, 118+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
 9, 18, 121+128, 
19, 28, 122+128, 
29, 38, 123+128, 
39, 48, 124+128, 
49, 58, 125+128, 
59, 69, 126+128, 
70, 80, 127+128, 
 8, 68, 79, 120+128, 
 0, 20, 40, 60, 104+128, 
10, 30, 50, 71, 105+128, 
 1, 21, 41, 61, 106+128, 
11, 31, 51, 72, 107+128, 
 2, 22, 42, 62, 108+128, 
12, 32, 52, 73, 109+128, 
 3, 23, 43, 63, 110+128, 
13, 33, 53, 74, 111+128, 
 4, 24, 44, 64, 112+128, 
14, 34, 54, 75, 113+128, 
 5, 25, 45, 65, 114+128, 
15, 35, 55, 76, 115+128, 
 6, 26, 46, 66, 116+128, 
16, 36, 56, 77, 117+128, 
 7, 27, 47, 67, 118+128, 
17, 37, 57, 78, 119+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
13, 26, 123+128, 
27, 40, 124+128, 
41, 55, 125+128, 
56, 69, 126+128, 
70, 84, 127+128, 
12, 54, 83, 122+128, 
 0, 14, 28, 42, 104+128, 
 1, 15, 43, 71, 105+128, 
 2, 16, 29, 72, 106+128, 
 3, 17, 44, 73, 107+128, 
30, 45, 57, 74, 108+128, 
18, 31, 46, 58, 109+128, 
19, 32, 47, 59, 110+128, 
 4, 33, 48, 60, 111+128, 
 5, 20, 61, 75, 112+128, 
34, 49, 62, 76, 113+128, 
 6, 50, 63, 77, 114+128, 
21, 51, 64, 78, 115+128, 
 7, 35, 65, 79, 116+128, 
 8, 22, 66, 80, 117+128, 
 9, 23, 36, 67, 118+128, 
10, 24, 37, 68, 119+128, 
25, 38, 52, 81, 120+128, 
11, 39, 53, 82, 121+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
13, 27, 123+128, 
28, 42, 124+128, 
43, 57, 125+128, 
58, 71, 126+128, 
72, 87, 127+128, 
14, 44, 73, 104+128, 
 0, 45, 59, 105+128, 
15, 29, 60, 106+128, 
 1, 16, 61, 107+128, 
17, 46, 74, 108+128, 
30, 62, 75, 109+128, 
 2, 31, 63, 110+128, 
 3, 47, 76, 111+128, 
 4, 32, 48, 112+128, 
18, 33, 77, 113+128, 
19, 49, 78, 114+128, 
12, 41, 86, 122+128, 
 5, 20, 34, 50, 64, 79, 115+128, 
 6, 21, 35, 51, 65, 80, 116+128, 
 7, 22, 36, 52, 66, 81, 117+128, 
 8, 23, 37, 53, 67, 82, 118+128, 
 9, 24, 38, 54, 68, 83, 119+128, 
10, 25, 39, 55, 69, 84, 120+128, 
11, 26, 40, 56, 70, 85, 121+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
19, 38, 125+128, 
39, 58, 126+128, 
59, 79, 127+128, 
 0, 40, 60, 104+128, 
 1, 20, 41, 105+128, 
 2, 42, 61, 106+128, 
21, 43, 62, 107+128, 
 3, 22, 44, 108+128, 
 4, 23, 63, 109+128, 
24, 45, 64, 110+128, 
 5, 25, 65, 111+128, 
 7, 47, 67, 113+128, 
18, 37, 78, 124+128, 
 6, 26, 46, 66, 112+128, 
 8, 27, 48, 68, 114+128, 
 9, 28, 49, 69, 115+128, 
10, 29, 50, 70, 116+128, 
11, 30, 51, 71, 117+128, 
12, 31, 52, 72, 118+128, 
13, 32, 53, 73, 119+128, 
14, 33, 54, 74, 120+128, 
15, 34, 55, 75, 121+128, 
16, 35, 56, 76, 122+128, 
17, 36, 57, 77, 123+128, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)) , 8 );
		end if;
	end process;
	
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity VNP_Output_Memory is
	generic(
		z			: integer := 96
	);
	Port (
		clk			: in  std_logic;
		
		RdAddr		: in  std_logic_vector(9 downto 0);
		Do			: out std_logic_vector(13 downto 0)
	);
end VNP_Output_Memory;

architecture Behavioral of VNP_Output_Memory is	
	------------------------------------O------------------------------------
	type ARRAY_TYPE is array (0 to 128*6-1) of integer;
	constant ROM 						: ARRAY_TYPE  := (
( 0*z/96)*128+ 5, ( 0*z/96)*128+11, ( 0*z/96)*128+117, 
( 0*z/96)*128+12, ( 0*z/96)*128+18, ( 0*z/96)*128+118, 
( 0*z/96)*128+19, ( 0*z/96)*128+24, ( 0*z/96)*128+119, 
( 0*z/96)*128+25, ( 0*z/96)*128+30, ( 0*z/96)*128+120, 
( 0*z/96)*128+31, ( 0*z/96)*128+37, ( 0*z/96)*128+121, 
( 0*z/96)*128+38, ( 0*z/96)*128+43, ( 0*z/96)*128+122, 
( 0*z/96)*128+44, ( 0*z/96)*128+49, ( 0*z/96)*128+123, 
( 0*z/96)*128+50, ( 0*z/96)*128+56, ( 0*z/96)*128+124, 
( 0*z/96)*128+57, ( 0*z/96)*128+62, ( 0*z/96)*128+125, 
( 0*z/96)*128+63, ( 0*z/96)*128+68, ( 0*z/96)*128+126, 
( 0*z/96)*128+69, ( 0*z/96)*128+75, ( 0*z/96)*128+127, 
(61*z/96)*128+20, (12*z/96)*128+51, (43*z/96)*128+70, ( 0*z/96)*128+104, 
(94*z/96)*128+ 0, (27*z/96)*128+ 6, (11*z/96)*128+45, ( 0*z/96)*128+105, 
(24*z/96)*128+13, (53*z/96)*128+40, (65*z/96)*128+65, ( 0*z/96)*128+107, 
(22*z/96)*128+14, (46*z/96)*128+32, (83*z/96)*128+52, ( 0*z/96)*128+108, 
(79*z/96)*128+ 8, (84*z/96)*128+27, ( 2*z/96)*128+47, ( 0*z/96)*128+110, 
(55*z/96)*128+ 2, (65*z/96)*128+22, (39*z/96)*128+66, ( 0*z/96)*128+112, 
(72*z/96)*128+29, (18*z/96)*128+42, (70*z/96)*128+60, ( 0*z/96)*128+114, 
( 7*z/96)*128+ 4, ( 0*z/96)*128+36, ( 7*z/96)*128+74, ( 0*z/96)*128+116, 
(73*z/96)*128+ 1, (47*z/96)*128+21, (39*z/96)*128+26, (95*z/96)*128+39, (73*z/96)*128+46, ( 7*z/96)*128+64, ( 0*z/96)*128+106, 
(22*z/96)*128+ 7, (81*z/96)*128+15, (40*z/96)*128+33, (24*z/96)*128+53, (94*z/96)*128+58, (66*z/96)*128+71, ( 0*z/96)*128+109, 
( 9*z/96)*128+ 9, (33*z/96)*128+16, (82*z/96)*128+34, (43*z/96)*128+54, (59*z/96)*128+59, (41*z/96)*128+72, ( 0*z/96)*128+111, 
(83*z/96)*128+ 3, (25*z/96)*128+23, (41*z/96)*128+28, (14*z/96)*128+41, (47*z/96)*128+48, (49*z/96)*128+67, ( 0*z/96)*128+113, 
(12*z/96)*128+10, ( 0*z/96)*128+17, (79*z/96)*128+35, (51*z/96)*128+55, (72*z/96)*128+61, (26*z/96)*128+73, ( 0*z/96)*128+115, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
( 0 mod z)*128+ 9, ( 0 mod z)*128+18, ( 0*z/96)*128+121, 
( 0 mod z)*128+19, ( 0 mod z)*128+28, ( 0*z/96)*128+122, 
( 0 mod z)*128+29, ( 0 mod z)*128+38, ( 0*z/96)*128+123, 
( 0 mod z)*128+39, ( 0 mod z)*128+48, ( 0*z/96)*128+124, 
( 0 mod z)*128+49, ( 0 mod z)*128+58, ( 0*z/96)*128+125, 
( 0 mod z)*128+59, ( 0 mod z)*128+68, ( 0*z/96)*128+126, 
( 0 mod z)*128+69, ( 0 mod z)*128+79, ( 0*z/96)*128+127, 
( 3 mod z)*128+ 0, (20 mod z)*128+40, (35 mod z)*128+60, ( 0*z/96)*128+104, 
( 0 mod z)*128+ 1, (25 mod z)*128+61, ( 6 mod z)*128+70, ( 0*z/96)*128+105, 
( 2 mod z)*128+21, (24 mod z)*128+31, (37 mod z)*128+62, ( 0*z/96)*128+107, 
( 2 mod z)*128+ 2, (36 mod z)*128+11, (28 mod z)*128+51, ( 0*z/96)*128+108, 
( 0 mod z)*128+33, (29 mod z)*128+43, ( 4 mod z)*128+72, ( 0*z/96)*128+110, 
( 3 mod z)*128+ 4, (34 mod z)*128+12, (40 mod z)*128+23, ( 0*z/96)*128+111, 
( 3 mod z)*128+24, (28 mod z)*128+44, (30 mod z)*128+74, ( 0*z/96)*128+113, 
( 1 mod z)*128+ 6, (17 mod z)*128+35, (36 mod z)*128+54, ( 0*z/96)*128+114, 
( 2 mod z)*128+15, ( 9 mod z)*128+55, (36 mod z)*128+76, ( 0*z/96)*128+116, 
( 2 mod z)*128+26, (38 mod z)*128+46, ( 4 mod z)*128+66, ( 0*z/96)*128+117, 
( 0 mod z)*128+17, (39 mod z)*128+37, (45 mod z)*128+57, ( 0*z/96)*128+119, 
( 1 mod z)*128+ 8, ( 0 mod z)*128+47, ( 1 mod z)*128+78, ( 0*z/96)*128+120, 
( 1 mod z)*128+10, (12 mod z)*128+20, (19 mod z)*128+30, ( 6 mod z)*128+41, (10 mod z)*128+50, ( 6 mod z)*128+71, ( 0*z/96)*128+106, 
( 0 mod z)*128+ 3, (15 mod z)*128+22, ( 3 mod z)*128+32, (10 mod z)*128+42, (20 mod z)*128+52, (21 mod z)*128+63, ( 0*z/96)*128+109, 
( 7 mod z)*128+ 5, (10 mod z)*128+13, ( 6 mod z)*128+34, ( 8 mod z)*128+53, ( 5 mod z)*128+64, (14 mod z)*128+73, ( 0*z/96)*128+112, 
( 1 mod z)*128+ 7, (18 mod z)*128+14, (15 mod z)*128+25, (14 mod z)*128+45, ( 0 mod z)*128+65, ( 3 mod z)*128+75, ( 0*z/96)*128+115, 
( 3 mod z)*128+16, (13 mod z)*128+27, ( 8 mod z)*128+36, (21 mod z)*128+56, (20 mod z)*128+67, (14 mod z)*128+77, ( 0*z/96)*128+118, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
( 0*z/96)*128+ 9, ( 0*z/96)*128+18, ( 0*z/96)*128+121, 
( 0*z/96)*128+19, ( 0*z/96)*128+28, ( 0*z/96)*128+122, 
( 0*z/96)*128+29, ( 0*z/96)*128+38, ( 0*z/96)*128+123, 
( 0*z/96)*128+39, ( 0*z/96)*128+48, ( 0*z/96)*128+124, 
( 0*z/96)*128+49, ( 0*z/96)*128+58, ( 0*z/96)*128+125, 
( 0*z/96)*128+59, ( 0*z/96)*128+69, ( 0*z/96)*128+126, 
( 0*z/96)*128+70, ( 0*z/96)*128+80, ( 0*z/96)*128+127, 
(95*z/96)*128+ 8, ( 0*z/96)*128+68, (95*z/96)*128+79, ( 0*z/96)*128+120, 
( 2*z/96)*128+ 0, (10*z/96)*128+20, (23*z/96)*128+40, (32*z/96)*128+60, ( 0*z/96)*128+104, 
(69*z/96)*128+10, (28*z/96)*128+30, (30*z/96)*128+50, ( 0*z/96)*128+71, ( 0*z/96)*128+105, 
(19*z/96)*128+ 1, (86*z/96)*128+21, (29*z/96)*128+41, ( 0*z/96)*128+61, ( 0*z/96)*128+106, 
(88*z/96)*128+11, (32*z/96)*128+31, (65*z/96)*128+51, (47*z/96)*128+72, ( 0*z/96)*128+107, 
(47*z/96)*128+ 2, (62*z/96)*128+22, (15*z/96)*128+42, (15*z/96)*128+62, ( 0*z/96)*128+108, 
(33*z/96)*128+12, (81*z/96)*128+32, (54*z/96)*128+52, (13*z/96)*128+73, ( 0*z/96)*128+109, 
(48*z/96)*128+ 3, (28*z/96)*128+23, (30*z/96)*128+43, (56*z/96)*128+63, ( 0*z/96)*128+110, 
( 3*z/96)*128+13, (27*z/96)*128+33, (14*z/96)*128+53, (61*z/96)*128+74, ( 0*z/96)*128+111, 
(36*z/96)*128+ 4, (85*z/96)*128+24, (66*z/96)*128+44, (85*z/96)*128+64, ( 0*z/96)*128+112, 
(16*z/96)*128+14, (88*z/96)*128+34, ( 0*z/96)*128+54, (84*z/96)*128+75, ( 0*z/96)*128+113, 
(82*z/96)*128+ 5, (16*z/96)*128+25, (24*z/96)*128+45, ( 5*z/96)*128+65, ( 0*z/96)*128+114, 
(37*z/96)*128+15, ( 5*z/96)*128+35, (30*z/96)*128+55, (55*z/96)*128+76, ( 0*z/96)*128+115, 
(47*z/96)*128+ 6, (34*z/96)*128+26, (50*z/96)*128+46, ( 6*z/96)*128+66, ( 0*z/96)*128+116, 
(40*z/96)*128+16, (56*z/96)*128+36, (74*z/96)*128+56, (78*z/96)*128+77, ( 0*z/96)*128+117, 
(15*z/96)*128+ 7, (73*z/96)*128+27, (62*z/96)*128+47, (52*z/96)*128+67, ( 0*z/96)*128+118, 
(48*z/96)*128+17, (37*z/96)*128+37, ( 0*z/96)*128+57, (41*z/96)*128+78, ( 0*z/96)*128+119, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
( 0*z/96)*128+13, ( 0*z/96)*128+26, ( 0*z/96)*128+123, 
( 0*z/96)*128+27, ( 0*z/96)*128+40, ( 0*z/96)*128+124, 
( 0*z/96)*128+41, ( 0*z/96)*128+55, ( 0*z/96)*128+125, 
( 0*z/96)*128+56, ( 0*z/96)*128+69, ( 0*z/96)*128+126, 
( 0*z/96)*128+70, ( 0*z/96)*128+84, ( 0*z/96)*128+127, 
(48*z/96)*128+12, ( 0*z/96)*128+54, (48*z/96)*128+83, ( 0*z/96)*128+122, 
( 6*z/96)*128+ 0, (62*z/96)*128+14, (71*z/96)*128+28, (38*z/96)*128+42, ( 0*z/96)*128+104, 
(38*z/96)*128+ 1, (94*z/96)*128+15, (61*z/96)*128+43, (63*z/96)*128+71, ( 0*z/96)*128+105, 
( 3*z/96)*128+ 2, (19*z/96)*128+16, (55*z/96)*128+29, (31*z/96)*128+72, ( 0*z/96)*128+106, 
(93*z/96)*128+ 3, (84*z/96)*128+17, (66*z/96)*128+44, (88*z/96)*128+73, ( 0*z/96)*128+107, 
(12*z/96)*128+30, ( 9*z/96)*128+45, (32*z/96)*128+57, (20*z/96)*128+74, ( 0*z/96)*128+108, 
(92*z/96)*128+18, (66*z/96)*128+31, (73*z/96)*128+46, (52*z/96)*128+58, ( 0*z/96)*128+109, 
(78*z/96)*128+19, (45*z/96)*128+32, (47*z/96)*128+47, (55*z/96)*128+59, ( 0*z/96)*128+110, 
(30*z/96)*128+ 4, (79*z/96)*128+33, (64*z/96)*128+48, (80*z/96)*128+60, ( 0*z/96)*128+111, 
(70*z/96)*128+ 5, (15*z/96)*128+20, (95*z/96)*128+61, ( 6*z/96)*128+75, ( 0*z/96)*128+112, 
(78*z/96)*128+34, (39*z/96)*128+49, (22*z/96)*128+62, (40*z/96)*128+76, ( 0*z/96)*128+113, 
(86*z/96)*128+ 6, (61*z/96)*128+50, ( 6*z/96)*128+63, (56*z/96)*128+77, ( 0*z/96)*128+114, 
(92*z/96)*128+21, (43*z/96)*128+51, (51*z/96)*128+64, (16*z/96)*128+78, ( 0*z/96)*128+115, 
(37*z/96)*128+ 7, (10*z/96)*128+35, (24*z/96)*128+65, (71*z/96)*128+79, ( 0*z/96)*128+116, 
(38*z/96)*128+ 8, (45*z/96)*128+22, (90*z/96)*128+66, (53*z/96)*128+80, ( 0*z/96)*128+117, 
( 4*z/96)*128+ 9, (24*z/96)*128+23, (22*z/96)*128+36, (44*z/96)*128+67, ( 0*z/96)*128+118, 
(11*z/96)*128+10, (32*z/96)*128+24, (55*z/96)*128+37, (20*z/96)*128+68, ( 0*z/96)*128+119, 
(30*z/96)*128+25, (70*z/96)*128+38, (95*z/96)*128+52, (27*z/96)*128+81, ( 0*z/96)*128+120, 
(46*z/96)*128+11, (82*z/96)*128+39, (32*z/96)*128+53, (26*z/96)*128+82, ( 0*z/96)*128+121, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
( 0*z/96)*128+13, ( 0*z/96)*128+27, ( 0*z/96)*128+123, 
( 0*z/96)*128+28, ( 0*z/96)*128+42, ( 0*z/96)*128+124, 
( 0*z/96)*128+43, ( 0*z/96)*128+57, ( 0*z/96)*128+125, 
( 0*z/96)*128+58, ( 0*z/96)*128+71, ( 0*z/96)*128+126, 
( 0*z/96)*128+72, ( 0*z/96)*128+87, ( 0*z/96)*128+127, 
(42*z/96)*128+14, (64*z/96)*128+44, (77*z/96)*128+73, ( 0*z/96)*128+104, 
(81*z/96)*128+ 0, ( 2*z/96)*128+45, (53*z/96)*128+59, ( 0*z/96)*128+105, 
(14*z/96)*128+15, (20*z/96)*128+29, (60*z/96)*128+60, ( 0*z/96)*128+106, 
(28*z/96)*128+ 1, (68*z/96)*128+16, (80*z/96)*128+61, ( 0*z/96)*128+107, 
(32*z/96)*128+17, (63*z/96)*128+46, (15*z/96)*128+74, ( 0*z/96)*128+108, 
(63*z/96)*128+30, (26*z/96)*128+62, (28*z/96)*128+75, ( 0*z/96)*128+109, 
(14*z/96)*128+ 2, (39*z/96)*128+31, (75*z/96)*128+63, ( 0*z/96)*128+110, 
(25*z/96)*128+ 3, ( 3*z/96)*128+47, (35*z/96)*128+76, ( 0*z/96)*128+111, 
(17*z/96)*128+ 4, (70*z/96)*128+32, (51*z/96)*128+48, ( 0*z/96)*128+112, 
(70*z/96)*128+18, (67*z/96)*128+33, (72*z/96)*128+77, ( 0*z/96)*128+113, 
(43*z/96)*128+19, (81*z/96)*128+49, (30*z/96)*128+78, ( 0*z/96)*128+114, 
( 0*z/96)*128+12, (80*z/96)*128+41, ( 0*z/96)*128+86, ( 0*z/96)*128+122, 
(85*z/96)*128+ 5, (11*z/96)*128+20, (38*z/96)*128+34, (15*z/96)*128+50, (86*z/96)*128+64, (68*z/96)*128+79, ( 0*z/96)*128+115, 
(29*z/96)*128+ 6, (36*z/96)*128+21, ( 4*z/96)*128+35, (94*z/96)*128+51, (77*z/96)*128+65, (85*z/96)*128+80, ( 0*z/96)*128+116, 
(52*z/96)*128+ 7, (40*z/96)*128+22, (72*z/96)*128+36, ( 9*z/96)*128+52, ( 1*z/96)*128+66, (84*z/96)*128+81, ( 0*z/96)*128+117, 
(78*z/96)*128+ 8, (33*z/96)*128+23, (47*z/96)*128+37, (85*z/96)*128+53, ( 3*z/96)*128+67, (26*z/96)*128+82, ( 0*z/96)*128+118, 
(95*z/96)*128+ 9, (57*z/96)*128+24, (29*z/96)*128+38, (36*z/96)*128+54, (72*z/96)*128+68, (64*z/96)*128+83, ( 0*z/96)*128+119, 
(22*z/96)*128+10, (38*z/96)*128+25, (60*z/96)*128+39, (14*z/96)*128+55, (60*z/96)*128+69, (11*z/96)*128+84, ( 0*z/96)*128+120, 
(92*z/96)*128+11, (24*z/96)*128+26, ( 5*z/96)*128+40, (19*z/96)*128+56, (25*z/96)*128+70, (89*z/96)*128+85, ( 0*z/96)*128+121, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
( 0*z/96)*128+19, ( 0*z/96)*128+38, ( 0*z/96)*128+125, 
( 0*z/96)*128+39, ( 0*z/96)*128+58, ( 0*z/96)*128+126, 
( 0*z/96)*128+59, ( 0*z/96)*128+79, ( 0*z/96)*128+127, 
( 1*z/96)*128+ 0, (51*z/96)*128+40, (50*z/96)*128+60, ( 0*z/96)*128+104, 
(25*z/96)*128+ 1, ( 6*z/96)*128+20, (81*z/96)*128+41, ( 0*z/96)*128+105, 
(55*z/96)*128+ 2, (83*z/96)*128+42, (50*z/96)*128+61, ( 0*z/96)*128+106, 
(36*z/96)*128+21, ( 4*z/96)*128+43, (15*z/96)*128+62, ( 0*z/96)*128+107, 
(47*z/96)*128+ 3, (40*z/96)*128+22, (67*z/96)*128+44, ( 0*z/96)*128+108, 
( 4*z/96)*128+ 4, (47*z/96)*128+23, (36*z/96)*128+63, ( 0*z/96)*128+109, 
(12*z/96)*128+24, (21*z/96)*128+45, (13*z/96)*128+64, ( 0*z/96)*128+110, 
(91*z/96)*128+ 5, (79*z/96)*128+25, (10*z/96)*128+65, ( 0*z/96)*128+111, 
( 8*z/96)*128+ 7, (24*z/96)*128+47, (20*z/96)*128+67, ( 0*z/96)*128+113, 
(80*z/96)*128+18, ( 0*z/96)*128+37, (80*z/96)*128+78, ( 0*z/96)*128+124, 
(84*z/96)*128+ 6, (47*z/96)*128+26, (31*z/96)*128+46, (11*z/96)*128+66, ( 0*z/96)*128+112, 
(86*z/96)*128+ 8, (41*z/96)*128+27, (91*z/96)*128+48, (53*z/96)*128+68, ( 0*z/96)*128+114, 
(52*z/96)*128+ 9, (21*z/96)*128+28, (61*z/96)*128+49, (90*z/96)*128+69, ( 0*z/96)*128+115, 
(82*z/96)*128+10, (12*z/96)*128+29, (81*z/96)*128+50, (29*z/96)*128+70, ( 0*z/96)*128+116, 
(33*z/96)*128+11, (71*z/96)*128+30, ( 9*z/96)*128+51, (92*z/96)*128+71, ( 0*z/96)*128+117, 
( 5*z/96)*128+12, (14*z/96)*128+31, (86*z/96)*128+52, (57*z/96)*128+72, ( 0*z/96)*128+118, 
( 0*z/96)*128+13, (72*z/96)*128+32, (78*z/96)*128+53, (30*z/96)*128+73, ( 0*z/96)*128+119, 
(36*z/96)*128+14, ( 0*z/96)*128+33, (60*z/96)*128+54, (84*z/96)*128+74, ( 0*z/96)*128+120, 
(20*z/96)*128+15, (44*z/96)*128+34, (88*z/96)*128+55, (92*z/96)*128+75, ( 0*z/96)*128+121, 
( 4*z/96)*128+16, (49*z/96)*128+35, (67*z/96)*128+56, (11*z/96)*128+76, ( 0*z/96)*128+122, 
(77*z/96)*128+17, ( 0*z/96)*128+36, (15*z/96)*128+57, (66*z/96)*128+77, ( 0*z/96)*128+123, 
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
);
begin
	process(clk)
	begin
		if rising_edge(clk) then
			Do <= conv_std_logic_vector( ROM(conv_integer(RdAddr)), 14);
		end if;
	end process;
	
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LLR_MEM is
	generic(
		z			: integer := 24;
		W			: integer := 8
	);
	Port (
		clk			: in  std_logic;

		WrDis		: in  std_logic;
		WrEn		: in  std_logic;
		WrAddr      : in  std_logic_vector(6 downto 0);
		Din         : in  std_logic_vector(z*W-1 downto 0);
		
		RdDis		: in  std_logic;
		RdEn		: in  std_logic;
		RdAddr      : in  std_logic_vector(6 downto 0);
		Dval		: out std_logic;
		Dout		: out std_logic_vector(z*W-1 downto 0)
	);
end LLR_MEM;

architecture Behavioral of LLR_MEM is
	------------------------------------O------------------------------------
	type fifo_type is array (0 to 127) of std_logic_vector(W*z-1 downto 0);
	signal fifo 						: fifo_type  := (others => (others => '0'));
	------------------------------------O------------------------------------
--	type ARRAY_TYPE_B is array (0 to z-1) of std_logic_vector(W-1 downto 0);
--	signal debug 						: ARRAY_TYPE_B  := (others => (others => '0'));
begin
--	-- synthesis translate_off
--	process(Din)
--	begin
--		for i in 0 to z-1 loop
--			debug(z-1-i) <= Din(W*(i+1)-1 downto W*i);
--		end loop;
--	end process;
--	-- synthesis translate_on
	process(clk)
	begin
		if rising_edge(clk) then
		    if WrEn = '1' then
				if WrDis = '0' or (WrDis = '1' and WrAddr < 104) then -- VNP'den gelen gereksiz yazma isteklerini engellemek icin, 104=128-24
					fifo(conv_integer(WrAddr)) <= Din;
				end if;
		    end if;
		
			Dval <= RdEn;
			Dout <= fifo(conv_integer(RdAddr));
			if RdDis = '1' and RdAddr < 104 then -- Ilk iterasyonda bellekte onceki pakete ait llr degerleri olacagi icin
				Dout <= (others => '0');
			end if;
		end if;
	end process;
	
end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity HD_MEM is
	generic(
		z						: integer := 96
	);
	Port (
		clk			: in  std_logic;

		WrEn		: in  std_logic;
		WrAddr      : in  std_logic_vector(6 downto 0);
		Din         : in  std_logic_vector(z-1 downto 0);

		RdEn		: in  std_logic;
		RdAddr      : in  std_logic_vector(6 downto 0);
		Dval		: out std_logic;
		Dout		: out std_logic_vector(z-1 downto 0)
	);
end HD_MEM;

architecture Behavioral of HD_MEM is
	------------------------------------O------------------------------------
	type fifo_type is array (0 to 127) of std_logic_vector(z-1 downto 0);
	signal fifo 						: fifo_type  := (others => (others => '0'));
	------------------------------------O------------------------------------
begin
	process(clk)
	begin
		if rising_edge(clk) then
		    if WrEn = '1' then
		        fifo(conv_integer(WrAddr)) <= Din;
		    end if;

			Dval <= RdEn;
			Dout <= fifo(conv_integer(RdAddr));
		end if;
	end process;

end Behavioral;
-------------------------------------------------------------------------------------
--=================================================================================--
--=================================================================================--
--=================================================================================--
-------------------------------------------------------------------------------------